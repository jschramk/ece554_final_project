module ExecuteMemoryPipe #() ();

endmodule