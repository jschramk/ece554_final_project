module PitchShift (
    input clk,
    input rst,
    input en,
    input [15:0]freq_domain_in[1023:0],
    output [15:0]freq_domain_out[1023:0],
    output ready_for_data,
    output done
);


endmodule