module FastFourierTransform (
    input clk,
    input rst,
    input [15:0]audio_in[2047:0],
    output [15:0]freq_domain_out[1023:0],
    output ready_for_data,
    output done
);


endmodule