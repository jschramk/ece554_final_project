module MemoryWritebackPipe #() ();

endmodule