module InverseFastFourierTransform (
    input clk,
    input rst,
    input [15:0]freq_domain_in[1023:0],
    output [15:0]audio_out[2047:0],
    output ready_for_data,
    output done
);


endmodule