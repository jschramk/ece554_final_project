module Memory #() ();

endmodule