module SineLUT (
    input [10:0] in, // mapping the sine function from [0, 2pi] to [0, 2047]
    output reg [15:0] out
);

always @(in) begin
    case(in)
        11'b00000000000 : out <= 16'sb00000000_00000000; // 0.00000
        11'b00000000001 : out <= 16'sb00000000_00000000; // 0.00307
        11'b00000000010 : out <= 16'sb00000000_00000001; // 0.00614
        11'b00000000011 : out <= 16'sb00000000_00000010; // 0.00920
        11'b00000000100 : out <= 16'sb00000000_00000011; // 0.01227
        11'b00000000101 : out <= 16'sb00000000_00000011; // 0.01534
        11'b00000000110 : out <= 16'sb00000000_00000100; // 0.01841
        11'b00000000111 : out <= 16'sb00000000_00000101; // 0.02147
        11'b00000001000 : out <= 16'sb00000000_00000110; // 0.02454
        11'b00000001001 : out <= 16'sb00000000_00000111; // 0.02761
        11'b00000001010 : out <= 16'sb00000000_00000111; // 0.03067
        11'b00000001011 : out <= 16'sb00000000_00001000; // 0.03374
        11'b00000001100 : out <= 16'sb00000000_00001001; // 0.03681
        11'b00000001101 : out <= 16'sb00000000_00001010; // 0.03987
        11'b00000001110 : out <= 16'sb00000000_00001010; // 0.04294
        11'b00000001111 : out <= 16'sb00000000_00001011; // 0.04600
        11'b00000010000 : out <= 16'sb00000000_00001100; // 0.04907
        11'b00000010001 : out <= 16'sb00000000_00001101; // 0.05213
        11'b00000010010 : out <= 16'sb00000000_00001110; // 0.05520
        11'b00000010011 : out <= 16'sb00000000_00001110; // 0.05826
        11'b00000010100 : out <= 16'sb00000000_00001111; // 0.06132
        11'b00000010101 : out <= 16'sb00000000_00010000; // 0.06438
        11'b00000010110 : out <= 16'sb00000000_00010001; // 0.06744
        11'b00000010111 : out <= 16'sb00000000_00010010; // 0.07050
        11'b00000011000 : out <= 16'sb00000000_00010010; // 0.07356
        11'b00000011001 : out <= 16'sb00000000_00010011; // 0.07662
        11'b00000011010 : out <= 16'sb00000000_00010100; // 0.07968
        11'b00000011011 : out <= 16'sb00000000_00010101; // 0.08274
        11'b00000011100 : out <= 16'sb00000000_00010101; // 0.08580
        11'b00000011101 : out <= 16'sb00000000_00010110; // 0.08885
        11'b00000011110 : out <= 16'sb00000000_00010111; // 0.09191
        11'b00000011111 : out <= 16'sb00000000_00011000; // 0.09496
        11'b00000100000 : out <= 16'sb00000000_00011001; // 0.09802
        11'b00000100001 : out <= 16'sb00000000_00011001; // 0.10107
        11'b00000100010 : out <= 16'sb00000000_00011010; // 0.10412
        11'b00000100011 : out <= 16'sb00000000_00011011; // 0.10717
        11'b00000100100 : out <= 16'sb00000000_00011100; // 0.11022
        11'b00000100101 : out <= 16'sb00000000_00011100; // 0.11327
        11'b00000100110 : out <= 16'sb00000000_00011101; // 0.11632
        11'b00000100111 : out <= 16'sb00000000_00011110; // 0.11937
        11'b00000101000 : out <= 16'sb00000000_00011111; // 0.12241
        11'b00000101001 : out <= 16'sb00000000_00100000; // 0.12545
        11'b00000101010 : out <= 16'sb00000000_00100000; // 0.12850
        11'b00000101011 : out <= 16'sb00000000_00100001; // 0.13154
        11'b00000101100 : out <= 16'sb00000000_00100010; // 0.13458
        11'b00000101101 : out <= 16'sb00000000_00100011; // 0.13762
        11'b00000101110 : out <= 16'sb00000000_00100100; // 0.14066
        11'b00000101111 : out <= 16'sb00000000_00100100; // 0.14370
        11'b00000110000 : out <= 16'sb00000000_00100101; // 0.14673
        11'b00000110001 : out <= 16'sb00000000_00100110; // 0.14976
        11'b00000110010 : out <= 16'sb00000000_00100111; // 0.15280
        11'b00000110011 : out <= 16'sb00000000_00100111; // 0.15583
        11'b00000110100 : out <= 16'sb00000000_00101000; // 0.15886
        11'b00000110101 : out <= 16'sb00000000_00101001; // 0.16189
        11'b00000110110 : out <= 16'sb00000000_00101010; // 0.16491
        11'b00000110111 : out <= 16'sb00000000_00101010; // 0.16794
        11'b00000111000 : out <= 16'sb00000000_00101011; // 0.17096
        11'b00000111001 : out <= 16'sb00000000_00101100; // 0.17398
        11'b00000111010 : out <= 16'sb00000000_00101101; // 0.17700
        11'b00000111011 : out <= 16'sb00000000_00101110; // 0.18002
        11'b00000111100 : out <= 16'sb00000000_00101110; // 0.18304
        11'b00000111101 : out <= 16'sb00000000_00101111; // 0.18606
        11'b00000111110 : out <= 16'sb00000000_00110000; // 0.18907
        11'b00000111111 : out <= 16'sb00000000_00110001; // 0.19208
        11'b00001000000 : out <= 16'sb00000000_00110001; // 0.19509
        11'b00001000001 : out <= 16'sb00000000_00110010; // 0.19810
        11'b00001000010 : out <= 16'sb00000000_00110011; // 0.20110
        11'b00001000011 : out <= 16'sb00000000_00110100; // 0.20411
        11'b00001000100 : out <= 16'sb00000000_00110101; // 0.20711
        11'b00001000101 : out <= 16'sb00000000_00110101; // 0.21011
        11'b00001000110 : out <= 16'sb00000000_00110110; // 0.21311
        11'b00001000111 : out <= 16'sb00000000_00110111; // 0.21611
        11'b00001001000 : out <= 16'sb00000000_00111000; // 0.21910
        11'b00001001001 : out <= 16'sb00000000_00111000; // 0.22209
        11'b00001001010 : out <= 16'sb00000000_00111001; // 0.22508
        11'b00001001011 : out <= 16'sb00000000_00111010; // 0.22807
        11'b00001001100 : out <= 16'sb00000000_00111011; // 0.23106
        11'b00001001101 : out <= 16'sb00000000_00111011; // 0.23404
        11'b00001001110 : out <= 16'sb00000000_00111100; // 0.23702
        11'b00001001111 : out <= 16'sb00000000_00111101; // 0.24000
        11'b00001010000 : out <= 16'sb00000000_00111110; // 0.24298
        11'b00001010001 : out <= 16'sb00000000_00111110; // 0.24596
        11'b00001010010 : out <= 16'sb00000000_00111111; // 0.24893
        11'b00001010011 : out <= 16'sb00000000_01000000; // 0.25190
        11'b00001010100 : out <= 16'sb00000000_01000001; // 0.25487
        11'b00001010101 : out <= 16'sb00000000_01000010; // 0.25783
        11'b00001010110 : out <= 16'sb00000000_01000010; // 0.26079
        11'b00001010111 : out <= 16'sb00000000_01000011; // 0.26375
        11'b00001011000 : out <= 16'sb00000000_01000100; // 0.26671
        11'b00001011001 : out <= 16'sb00000000_01000101; // 0.26967
        11'b00001011010 : out <= 16'sb00000000_01000101; // 0.27262
        11'b00001011011 : out <= 16'sb00000000_01000110; // 0.27557
        11'b00001011100 : out <= 16'sb00000000_01000111; // 0.27852
        11'b00001011101 : out <= 16'sb00000000_01001000; // 0.28146
        11'b00001011110 : out <= 16'sb00000000_01001000; // 0.28441
        11'b00001011111 : out <= 16'sb00000000_01001001; // 0.28735
        11'b00001100000 : out <= 16'sb00000000_01001010; // 0.29028
        11'b00001100001 : out <= 16'sb00000000_01001011; // 0.29322
        11'b00001100010 : out <= 16'sb00000000_01001011; // 0.29615
        11'b00001100011 : out <= 16'sb00000000_01001100; // 0.29908
        11'b00001100100 : out <= 16'sb00000000_01001101; // 0.30201
        11'b00001100101 : out <= 16'sb00000000_01001110; // 0.30493
        11'b00001100110 : out <= 16'sb00000000_01001110; // 0.30785
        11'b00001100111 : out <= 16'sb00000000_01001111; // 0.31077
        11'b00001101000 : out <= 16'sb00000000_01010000; // 0.31368
        11'b00001101001 : out <= 16'sb00000000_01010001; // 0.31659
        11'b00001101010 : out <= 16'sb00000000_01010001; // 0.31950
        11'b00001101011 : out <= 16'sb00000000_01010010; // 0.32241
        11'b00001101100 : out <= 16'sb00000000_01010011; // 0.32531
        11'b00001101101 : out <= 16'sb00000000_01010100; // 0.32821
        11'b00001101110 : out <= 16'sb00000000_01010100; // 0.33111
        11'b00001101111 : out <= 16'sb00000000_01010101; // 0.33400
        11'b00001110000 : out <= 16'sb00000000_01010110; // 0.33689
        11'b00001110001 : out <= 16'sb00000000_01010110; // 0.33978
        11'b00001110010 : out <= 16'sb00000000_01010111; // 0.34266
        11'b00001110011 : out <= 16'sb00000000_01011000; // 0.34554
        11'b00001110100 : out <= 16'sb00000000_01011001; // 0.34842
        11'b00001110101 : out <= 16'sb00000000_01011001; // 0.35129
        11'b00001110110 : out <= 16'sb00000000_01011010; // 0.35416
        11'b00001110111 : out <= 16'sb00000000_01011011; // 0.35703
        11'b00001111000 : out <= 16'sb00000000_01011100; // 0.35990
        11'b00001111001 : out <= 16'sb00000000_01011100; // 0.36276
        11'b00001111010 : out <= 16'sb00000000_01011101; // 0.36561
        11'b00001111011 : out <= 16'sb00000000_01011110; // 0.36847
        11'b00001111100 : out <= 16'sb00000000_01011111; // 0.37132
        11'b00001111101 : out <= 16'sb00000000_01011111; // 0.37416
        11'b00001111110 : out <= 16'sb00000000_01100000; // 0.37701
        11'b00001111111 : out <= 16'sb00000000_01100001; // 0.37985
        11'b00010000000 : out <= 16'sb00000000_01100001; // 0.38268
        11'b00010000001 : out <= 16'sb00000000_01100010; // 0.38552
        11'b00010000010 : out <= 16'sb00000000_01100011; // 0.38835
        11'b00010000011 : out <= 16'sb00000000_01100100; // 0.39117
        11'b00010000100 : out <= 16'sb00000000_01100100; // 0.39399
        11'b00010000101 : out <= 16'sb00000000_01100101; // 0.39681
        11'b00010000110 : out <= 16'sb00000000_01100110; // 0.39962
        11'b00010000111 : out <= 16'sb00000000_01100111; // 0.40243
        11'b00010001000 : out <= 16'sb00000000_01100111; // 0.40524
        11'b00010001001 : out <= 16'sb00000000_01101000; // 0.40804
        11'b00010001010 : out <= 16'sb00000000_01101001; // 0.41084
        11'b00010001011 : out <= 16'sb00000000_01101001; // 0.41364
        11'b00010001100 : out <= 16'sb00000000_01101010; // 0.41643
        11'b00010001101 : out <= 16'sb00000000_01101011; // 0.41922
        11'b00010001110 : out <= 16'sb00000000_01101100; // 0.42200
        11'b00010001111 : out <= 16'sb00000000_01101100; // 0.42478
        11'b00010010000 : out <= 16'sb00000000_01101101; // 0.42756
        11'b00010010001 : out <= 16'sb00000000_01101110; // 0.43033
        11'b00010010010 : out <= 16'sb00000000_01101110; // 0.43309
        11'b00010010011 : out <= 16'sb00000000_01101111; // 0.43586
        11'b00010010100 : out <= 16'sb00000000_01110000; // 0.43862
        11'b00010010101 : out <= 16'sb00000000_01110000; // 0.44137
        11'b00010010110 : out <= 16'sb00000000_01110001; // 0.44412
        11'b00010010111 : out <= 16'sb00000000_01110010; // 0.44687
        11'b00010011000 : out <= 16'sb00000000_01110011; // 0.44961
        11'b00010011001 : out <= 16'sb00000000_01110011; // 0.45235
        11'b00010011010 : out <= 16'sb00000000_01110100; // 0.45508
        11'b00010011011 : out <= 16'sb00000000_01110101; // 0.45781
        11'b00010011100 : out <= 16'sb00000000_01110101; // 0.46054
        11'b00010011101 : out <= 16'sb00000000_01110110; // 0.46326
        11'b00010011110 : out <= 16'sb00000000_01110111; // 0.46598
        11'b00010011111 : out <= 16'sb00000000_01110111; // 0.46869
        11'b00010100000 : out <= 16'sb00000000_01111000; // 0.47140
        11'b00010100001 : out <= 16'sb00000000_01111001; // 0.47410
        11'b00010100010 : out <= 16'sb00000000_01111010; // 0.47680
        11'b00010100011 : out <= 16'sb00000000_01111010; // 0.47949
        11'b00010100100 : out <= 16'sb00000000_01111011; // 0.48218
        11'b00010100101 : out <= 16'sb00000000_01111100; // 0.48487
        11'b00010100110 : out <= 16'sb00000000_01111100; // 0.48755
        11'b00010100111 : out <= 16'sb00000000_01111101; // 0.49023
        11'b00010101000 : out <= 16'sb00000000_01111110; // 0.49290
        11'b00010101001 : out <= 16'sb00000000_01111110; // 0.49557
        11'b00010101010 : out <= 16'sb00000000_01111111; // 0.49823
        11'b00010101011 : out <= 16'sb00000000_10000000; // 0.50089
        11'b00010101100 : out <= 16'sb00000000_10000000; // 0.50354
        11'b00010101101 : out <= 16'sb00000000_10000001; // 0.50619
        11'b00010101110 : out <= 16'sb00000000_10000010; // 0.50883
        11'b00010101111 : out <= 16'sb00000000_10000010; // 0.51147
        11'b00010110000 : out <= 16'sb00000000_10000011; // 0.51410
        11'b00010110001 : out <= 16'sb00000000_10000100; // 0.51673
        11'b00010110010 : out <= 16'sb00000000_10000100; // 0.51936
        11'b00010110011 : out <= 16'sb00000000_10000101; // 0.52198
        11'b00010110100 : out <= 16'sb00000000_10000110; // 0.52459
        11'b00010110101 : out <= 16'sb00000000_10000110; // 0.52720
        11'b00010110110 : out <= 16'sb00000000_10000111; // 0.52980
        11'b00010110111 : out <= 16'sb00000000_10001000; // 0.53240
        11'b00010111000 : out <= 16'sb00000000_10001000; // 0.53500
        11'b00010111001 : out <= 16'sb00000000_10001001; // 0.53759
        11'b00010111010 : out <= 16'sb00000000_10001010; // 0.54017
        11'b00010111011 : out <= 16'sb00000000_10001010; // 0.54275
        11'b00010111100 : out <= 16'sb00000000_10001011; // 0.54532
        11'b00010111101 : out <= 16'sb00000000_10001100; // 0.54789
        11'b00010111110 : out <= 16'sb00000000_10001100; // 0.55046
        11'b00010111111 : out <= 16'sb00000000_10001101; // 0.55302
        11'b00011000000 : out <= 16'sb00000000_10001110; // 0.55557
        11'b00011000001 : out <= 16'sb00000000_10001110; // 0.55812
        11'b00011000010 : out <= 16'sb00000000_10001111; // 0.56066
        11'b00011000011 : out <= 16'sb00000000_10010000; // 0.56320
        11'b00011000100 : out <= 16'sb00000000_10010000; // 0.56573
        11'b00011000101 : out <= 16'sb00000000_10010001; // 0.56826
        11'b00011000110 : out <= 16'sb00000000_10010010; // 0.57078
        11'b00011000111 : out <= 16'sb00000000_10010010; // 0.57330
        11'b00011001000 : out <= 16'sb00000000_10010011; // 0.57581
        11'b00011001001 : out <= 16'sb00000000_10010100; // 0.57831
        11'b00011001010 : out <= 16'sb00000000_10010100; // 0.58081
        11'b00011001011 : out <= 16'sb00000000_10010101; // 0.58331
        11'b00011001100 : out <= 16'sb00000000_10010101; // 0.58580
        11'b00011001101 : out <= 16'sb00000000_10010110; // 0.58828
        11'b00011001110 : out <= 16'sb00000000_10010111; // 0.59076
        11'b00011001111 : out <= 16'sb00000000_10010111; // 0.59323
        11'b00011010000 : out <= 16'sb00000000_10011000; // 0.59570
        11'b00011010001 : out <= 16'sb00000000_10011001; // 0.59816
        11'b00011010010 : out <= 16'sb00000000_10011001; // 0.60062
        11'b00011010011 : out <= 16'sb00000000_10011010; // 0.60307
        11'b00011010100 : out <= 16'sb00000000_10011011; // 0.60551
        11'b00011010101 : out <= 16'sb00000000_10011011; // 0.60795
        11'b00011010110 : out <= 16'sb00000000_10011100; // 0.61038
        11'b00011010111 : out <= 16'sb00000000_10011100; // 0.61281
        11'b00011011000 : out <= 16'sb00000000_10011101; // 0.61523
        11'b00011011001 : out <= 16'sb00000000_10011110; // 0.61765
        11'b00011011010 : out <= 16'sb00000000_10011110; // 0.62006
        11'b00011011011 : out <= 16'sb00000000_10011111; // 0.62246
        11'b00011011100 : out <= 16'sb00000000_10011111; // 0.62486
        11'b00011011101 : out <= 16'sb00000000_10100000; // 0.62725
        11'b00011011110 : out <= 16'sb00000000_10100001; // 0.62964
        11'b00011011111 : out <= 16'sb00000000_10100001; // 0.63202
        11'b00011100000 : out <= 16'sb00000000_10100010; // 0.63439
        11'b00011100001 : out <= 16'sb00000000_10100011; // 0.63676
        11'b00011100010 : out <= 16'sb00000000_10100011; // 0.63912
        11'b00011100011 : out <= 16'sb00000000_10100100; // 0.64148
        11'b00011100100 : out <= 16'sb00000000_10100100; // 0.64383
        11'b00011100101 : out <= 16'sb00000000_10100101; // 0.64618
        11'b00011100110 : out <= 16'sb00000000_10100110; // 0.64851
        11'b00011100111 : out <= 16'sb00000000_10100110; // 0.65085
        11'b00011101000 : out <= 16'sb00000000_10100111; // 0.65317
        11'b00011101001 : out <= 16'sb00000000_10100111; // 0.65549
        11'b00011101010 : out <= 16'sb00000000_10101000; // 0.65781
        11'b00011101011 : out <= 16'sb00000000_10101000; // 0.66011
        11'b00011101100 : out <= 16'sb00000000_10101001; // 0.66242
        11'b00011101101 : out <= 16'sb00000000_10101010; // 0.66471
        11'b00011101110 : out <= 16'sb00000000_10101010; // 0.66700
        11'b00011101111 : out <= 16'sb00000000_10101011; // 0.66928
        11'b00011110000 : out <= 16'sb00000000_10101011; // 0.67156
        11'b00011110001 : out <= 16'sb00000000_10101100; // 0.67383
        11'b00011110010 : out <= 16'sb00000000_10101101; // 0.67609
        11'b00011110011 : out <= 16'sb00000000_10101101; // 0.67835
        11'b00011110100 : out <= 16'sb00000000_10101110; // 0.68060
        11'b00011110101 : out <= 16'sb00000000_10101110; // 0.68285
        11'b00011110110 : out <= 16'sb00000000_10101111; // 0.68508
        11'b00011110111 : out <= 16'sb00000000_10101111; // 0.68732
        11'b00011111000 : out <= 16'sb00000000_10110000; // 0.68954
        11'b00011111001 : out <= 16'sb00000000_10110001; // 0.69176
        11'b00011111010 : out <= 16'sb00000000_10110001; // 0.69397
        11'b00011111011 : out <= 16'sb00000000_10110010; // 0.69618
        11'b00011111100 : out <= 16'sb00000000_10110010; // 0.69838
        11'b00011111101 : out <= 16'sb00000000_10110011; // 0.70057
        11'b00011111110 : out <= 16'sb00000000_10110011; // 0.70275
        11'b00011111111 : out <= 16'sb00000000_10110100; // 0.70493
        11'b00100000000 : out <= 16'sb00000000_10110101; // 0.70711
        11'b00100000001 : out <= 16'sb00000000_10110101; // 0.70927
        11'b00100000010 : out <= 16'sb00000000_10110110; // 0.71143
        11'b00100000011 : out <= 16'sb00000000_10110110; // 0.71358
        11'b00100000100 : out <= 16'sb00000000_10110111; // 0.71573
        11'b00100000101 : out <= 16'sb00000000_10110111; // 0.71787
        11'b00100000110 : out <= 16'sb00000000_10111000; // 0.72000
        11'b00100000111 : out <= 16'sb00000000_10111000; // 0.72213
        11'b00100001000 : out <= 16'sb00000000_10111001; // 0.72425
        11'b00100001001 : out <= 16'sb00000000_10111001; // 0.72636
        11'b00100001010 : out <= 16'sb00000000_10111010; // 0.72846
        11'b00100001011 : out <= 16'sb00000000_10111011; // 0.73056
        11'b00100001100 : out <= 16'sb00000000_10111011; // 0.73265
        11'b00100001101 : out <= 16'sb00000000_10111100; // 0.73474
        11'b00100001110 : out <= 16'sb00000000_10111100; // 0.73682
        11'b00100001111 : out <= 16'sb00000000_10111101; // 0.73889
        11'b00100010000 : out <= 16'sb00000000_10111101; // 0.74095
        11'b00100010001 : out <= 16'sb00000000_10111110; // 0.74301
        11'b00100010010 : out <= 16'sb00000000_10111110; // 0.74506
        11'b00100010011 : out <= 16'sb00000000_10111111; // 0.74710
        11'b00100010100 : out <= 16'sb00000000_10111111; // 0.74914
        11'b00100010101 : out <= 16'sb00000000_11000000; // 0.75117
        11'b00100010110 : out <= 16'sb00000000_11000000; // 0.75319
        11'b00100010111 : out <= 16'sb00000000_11000001; // 0.75520
        11'b00100011000 : out <= 16'sb00000000_11000001; // 0.75721
        11'b00100011001 : out <= 16'sb00000000_11000010; // 0.75921
        11'b00100011010 : out <= 16'sb00000000_11000010; // 0.76120
        11'b00100011011 : out <= 16'sb00000000_11000011; // 0.76319
        11'b00100011100 : out <= 16'sb00000000_11000011; // 0.76517
        11'b00100011101 : out <= 16'sb00000000_11000100; // 0.76714
        11'b00100011110 : out <= 16'sb00000000_11000100; // 0.76910
        11'b00100011111 : out <= 16'sb00000000_11000101; // 0.77106
        11'b00100100000 : out <= 16'sb00000000_11000101; // 0.77301
        11'b00100100001 : out <= 16'sb00000000_11000110; // 0.77495
        11'b00100100010 : out <= 16'sb00000000_11000110; // 0.77689
        11'b00100100011 : out <= 16'sb00000000_11000111; // 0.77882
        11'b00100100100 : out <= 16'sb00000000_11000111; // 0.78074
        11'b00100100101 : out <= 16'sb00000000_11001000; // 0.78265
        11'b00100100110 : out <= 16'sb00000000_11001000; // 0.78456
        11'b00100100111 : out <= 16'sb00000000_11001001; // 0.78646
        11'b00100101000 : out <= 16'sb00000000_11001001; // 0.78835
        11'b00100101001 : out <= 16'sb00000000_11001010; // 0.79023
        11'b00100101010 : out <= 16'sb00000000_11001010; // 0.79211
        11'b00100101011 : out <= 16'sb00000000_11001011; // 0.79398
        11'b00100101100 : out <= 16'sb00000000_11001011; // 0.79584
        11'b00100101101 : out <= 16'sb00000000_11001100; // 0.79769
        11'b00100101110 : out <= 16'sb00000000_11001100; // 0.79954
        11'b00100101111 : out <= 16'sb00000000_11001101; // 0.80138
        11'b00100110000 : out <= 16'sb00000000_11001101; // 0.80321
        11'b00100110001 : out <= 16'sb00000000_11001110; // 0.80503
        11'b00100110010 : out <= 16'sb00000000_11001110; // 0.80685
        11'b00100110011 : out <= 16'sb00000000_11001111; // 0.80866
        11'b00100110100 : out <= 16'sb00000000_11001111; // 0.81046
        11'b00100110101 : out <= 16'sb00000000_11001111; // 0.81225
        11'b00100110110 : out <= 16'sb00000000_11010000; // 0.81404
        11'b00100110111 : out <= 16'sb00000000_11010000; // 0.81581
        11'b00100111000 : out <= 16'sb00000000_11010001; // 0.81758
        11'b00100111001 : out <= 16'sb00000000_11010001; // 0.81935
        11'b00100111010 : out <= 16'sb00000000_11010010; // 0.82110
        11'b00100111011 : out <= 16'sb00000000_11010010; // 0.82285
        11'b00100111100 : out <= 16'sb00000000_11010011; // 0.82459
        11'b00100111101 : out <= 16'sb00000000_11010011; // 0.82632
        11'b00100111110 : out <= 16'sb00000000_11010011; // 0.82805
        11'b00100111111 : out <= 16'sb00000000_11010100; // 0.82976
        11'b00101000000 : out <= 16'sb00000000_11010100; // 0.83147
        11'b00101000001 : out <= 16'sb00000000_11010101; // 0.83317
        11'b00101000010 : out <= 16'sb00000000_11010101; // 0.83486
        11'b00101000011 : out <= 16'sb00000000_11010110; // 0.83655
        11'b00101000100 : out <= 16'sb00000000_11010110; // 0.83822
        11'b00101000101 : out <= 16'sb00000000_11010111; // 0.83989
        11'b00101000110 : out <= 16'sb00000000_11010111; // 0.84155
        11'b00101000111 : out <= 16'sb00000000_11010111; // 0.84321
        11'b00101001000 : out <= 16'sb00000000_11011000; // 0.84485
        11'b00101001001 : out <= 16'sb00000000_11011000; // 0.84649
        11'b00101001010 : out <= 16'sb00000000_11011001; // 0.84812
        11'b00101001011 : out <= 16'sb00000000_11011001; // 0.84974
        11'b00101001100 : out <= 16'sb00000000_11011001; // 0.85136
        11'b00101001101 : out <= 16'sb00000000_11011010; // 0.85296
        11'b00101001110 : out <= 16'sb00000000_11011010; // 0.85456
        11'b00101001111 : out <= 16'sb00000000_11011011; // 0.85615
        11'b00101010000 : out <= 16'sb00000000_11011011; // 0.85773
        11'b00101010001 : out <= 16'sb00000000_11011011; // 0.85930
        11'b00101010010 : out <= 16'sb00000000_11011100; // 0.86087
        11'b00101010011 : out <= 16'sb00000000_11011100; // 0.86242
        11'b00101010100 : out <= 16'sb00000000_11011101; // 0.86397
        11'b00101010101 : out <= 16'sb00000000_11011101; // 0.86551
        11'b00101010110 : out <= 16'sb00000000_11011101; // 0.86705
        11'b00101010111 : out <= 16'sb00000000_11011110; // 0.86857
        11'b00101011000 : out <= 16'sb00000000_11011110; // 0.87009
        11'b00101011001 : out <= 16'sb00000000_11011111; // 0.87160
        11'b00101011010 : out <= 16'sb00000000_11011111; // 0.87309
        11'b00101011011 : out <= 16'sb00000000_11011111; // 0.87459
        11'b00101011100 : out <= 16'sb00000000_11100000; // 0.87607
        11'b00101011101 : out <= 16'sb00000000_11100000; // 0.87755
        11'b00101011110 : out <= 16'sb00000000_11100001; // 0.87901
        11'b00101011111 : out <= 16'sb00000000_11100001; // 0.88047
        11'b00101100000 : out <= 16'sb00000000_11100001; // 0.88192
        11'b00101100001 : out <= 16'sb00000000_11100010; // 0.88336
        11'b00101100010 : out <= 16'sb00000000_11100010; // 0.88480
        11'b00101100011 : out <= 16'sb00000000_11100010; // 0.88622
        11'b00101100100 : out <= 16'sb00000000_11100011; // 0.88764
        11'b00101100101 : out <= 16'sb00000000_11100011; // 0.88905
        11'b00101100110 : out <= 16'sb00000000_11100011; // 0.89045
        11'b00101100111 : out <= 16'sb00000000_11100100; // 0.89184
        11'b00101101000 : out <= 16'sb00000000_11100100; // 0.89322
        11'b00101101001 : out <= 16'sb00000000_11100101; // 0.89460
        11'b00101101010 : out <= 16'sb00000000_11100101; // 0.89597
        11'b00101101011 : out <= 16'sb00000000_11100101; // 0.89732
        11'b00101101100 : out <= 16'sb00000000_11100110; // 0.89867
        11'b00101101101 : out <= 16'sb00000000_11100110; // 0.90002
        11'b00101101110 : out <= 16'sb00000000_11100110; // 0.90135
        11'b00101101111 : out <= 16'sb00000000_11100111; // 0.90267
        11'b00101110000 : out <= 16'sb00000000_11100111; // 0.90399
        11'b00101110001 : out <= 16'sb00000000_11100111; // 0.90530
        11'b00101110010 : out <= 16'sb00000000_11101000; // 0.90660
        11'b00101110011 : out <= 16'sb00000000_11101000; // 0.90789
        11'b00101110100 : out <= 16'sb00000000_11101000; // 0.90917
        11'b00101110101 : out <= 16'sb00000000_11101001; // 0.91044
        11'b00101110110 : out <= 16'sb00000000_11101001; // 0.91171
        11'b00101110111 : out <= 16'sb00000000_11101001; // 0.91296
        11'b00101111000 : out <= 16'sb00000000_11101010; // 0.91421
        11'b00101111001 : out <= 16'sb00000000_11101010; // 0.91545
        11'b00101111010 : out <= 16'sb00000000_11101010; // 0.91668
        11'b00101111011 : out <= 16'sb00000000_11101010; // 0.91790
        11'b00101111100 : out <= 16'sb00000000_11101011; // 0.91911
        11'b00101111101 : out <= 16'sb00000000_11101011; // 0.92032
        11'b00101111110 : out <= 16'sb00000000_11101011; // 0.92151
        11'b00101111111 : out <= 16'sb00000000_11101100; // 0.92270
        11'b00110000000 : out <= 16'sb00000000_11101100; // 0.92388
        11'b00110000001 : out <= 16'sb00000000_11101100; // 0.92505
        11'b00110000010 : out <= 16'sb00000000_11101101; // 0.92621
        11'b00110000011 : out <= 16'sb00000000_11101101; // 0.92736
        11'b00110000100 : out <= 16'sb00000000_11101101; // 0.92851
        11'b00110000101 : out <= 16'sb00000000_11101101; // 0.92964
        11'b00110000110 : out <= 16'sb00000000_11101110; // 0.93077
        11'b00110000111 : out <= 16'sb00000000_11101110; // 0.93188
        11'b00110001000 : out <= 16'sb00000000_11101110; // 0.93299
        11'b00110001001 : out <= 16'sb00000000_11101111; // 0.93409
        11'b00110001010 : out <= 16'sb00000000_11101111; // 0.93518
        11'b00110001011 : out <= 16'sb00000000_11101111; // 0.93627
        11'b00110001100 : out <= 16'sb00000000_11101111; // 0.93734
        11'b00110001101 : out <= 16'sb00000000_11110000; // 0.93840
        11'b00110001110 : out <= 16'sb00000000_11110000; // 0.93946
        11'b00110001111 : out <= 16'sb00000000_11110000; // 0.94051
        11'b00110010000 : out <= 16'sb00000000_11110001; // 0.94154
        11'b00110010001 : out <= 16'sb00000000_11110001; // 0.94257
        11'b00110010010 : out <= 16'sb00000000_11110001; // 0.94359
        11'b00110010011 : out <= 16'sb00000000_11110001; // 0.94460
        11'b00110010100 : out <= 16'sb00000000_11110010; // 0.94561
        11'b00110010101 : out <= 16'sb00000000_11110010; // 0.94660
        11'b00110010110 : out <= 16'sb00000000_11110010; // 0.94759
        11'b00110010111 : out <= 16'sb00000000_11110010; // 0.94856
        11'b00110011000 : out <= 16'sb00000000_11110011; // 0.94953
        11'b00110011001 : out <= 16'sb00000000_11110011; // 0.95049
        11'b00110011010 : out <= 16'sb00000000_11110011; // 0.95144
        11'b00110011011 : out <= 16'sb00000000_11110011; // 0.95238
        11'b00110011100 : out <= 16'sb00000000_11110100; // 0.95331
        11'b00110011101 : out <= 16'sb00000000_11110100; // 0.95423
        11'b00110011110 : out <= 16'sb00000000_11110100; // 0.95514
        11'b00110011111 : out <= 16'sb00000000_11110100; // 0.95605
        11'b00110100000 : out <= 16'sb00000000_11110100; // 0.95694
        11'b00110100001 : out <= 16'sb00000000_11110101; // 0.95783
        11'b00110100010 : out <= 16'sb00000000_11110101; // 0.95870
        11'b00110100011 : out <= 16'sb00000000_11110101; // 0.95957
        11'b00110100100 : out <= 16'sb00000000_11110101; // 0.96043
        11'b00110100101 : out <= 16'sb00000000_11110110; // 0.96128
        11'b00110100110 : out <= 16'sb00000000_11110110; // 0.96212
        11'b00110100111 : out <= 16'sb00000000_11110110; // 0.96295
        11'b00110101000 : out <= 16'sb00000000_11110110; // 0.96378
        11'b00110101001 : out <= 16'sb00000000_11110110; // 0.96459
        11'b00110101010 : out <= 16'sb00000000_11110111; // 0.96539
        11'b00110101011 : out <= 16'sb00000000_11110111; // 0.96619
        11'b00110101100 : out <= 16'sb00000000_11110111; // 0.96698
        11'b00110101101 : out <= 16'sb00000000_11110111; // 0.96775
        11'b00110101110 : out <= 16'sb00000000_11110111; // 0.96852
        11'b00110101111 : out <= 16'sb00000000_11111000; // 0.96928
        11'b00110110000 : out <= 16'sb00000000_11111000; // 0.97003
        11'b00110110001 : out <= 16'sb00000000_11111000; // 0.97077
        11'b00110110010 : out <= 16'sb00000000_11111000; // 0.97150
        11'b00110110011 : out <= 16'sb00000000_11111000; // 0.97223
        11'b00110110100 : out <= 16'sb00000000_11111001; // 0.97294
        11'b00110110101 : out <= 16'sb00000000_11111001; // 0.97364
        11'b00110110110 : out <= 16'sb00000000_11111001; // 0.97434
        11'b00110110111 : out <= 16'sb00000000_11111001; // 0.97503
        11'b00110111000 : out <= 16'sb00000000_11111001; // 0.97570
        11'b00110111001 : out <= 16'sb00000000_11111001; // 0.97637
        11'b00110111010 : out <= 16'sb00000000_11111010; // 0.97703
        11'b00110111011 : out <= 16'sb00000000_11111010; // 0.97768
        11'b00110111100 : out <= 16'sb00000000_11111010; // 0.97832
        11'b00110111101 : out <= 16'sb00000000_11111010; // 0.97895
        11'b00110111110 : out <= 16'sb00000000_11111010; // 0.97957
        11'b00110111111 : out <= 16'sb00000000_11111010; // 0.98018
        11'b00111000000 : out <= 16'sb00000000_11111011; // 0.98079
        11'b00111000001 : out <= 16'sb00000000_11111011; // 0.98138
        11'b00111000010 : out <= 16'sb00000000_11111011; // 0.98196
        11'b00111000011 : out <= 16'sb00000000_11111011; // 0.98254
        11'b00111000100 : out <= 16'sb00000000_11111011; // 0.98311
        11'b00111000101 : out <= 16'sb00000000_11111011; // 0.98366
        11'b00111000110 : out <= 16'sb00000000_11111011; // 0.98421
        11'b00111000111 : out <= 16'sb00000000_11111100; // 0.98475
        11'b00111001000 : out <= 16'sb00000000_11111100; // 0.98528
        11'b00111001001 : out <= 16'sb00000000_11111100; // 0.98580
        11'b00111001010 : out <= 16'sb00000000_11111100; // 0.98631
        11'b00111001011 : out <= 16'sb00000000_11111100; // 0.98681
        11'b00111001100 : out <= 16'sb00000000_11111100; // 0.98730
        11'b00111001101 : out <= 16'sb00000000_11111100; // 0.98778
        11'b00111001110 : out <= 16'sb00000000_11111100; // 0.98826
        11'b00111001111 : out <= 16'sb00000000_11111101; // 0.98872
        11'b00111010000 : out <= 16'sb00000000_11111101; // 0.98918
        11'b00111010001 : out <= 16'sb00000000_11111101; // 0.98962
        11'b00111010010 : out <= 16'sb00000000_11111101; // 0.99006
        11'b00111010011 : out <= 16'sb00000000_11111101; // 0.99049
        11'b00111010100 : out <= 16'sb00000000_11111101; // 0.99090
        11'b00111010101 : out <= 16'sb00000000_11111101; // 0.99131
        11'b00111010110 : out <= 16'sb00000000_11111101; // 0.99171
        11'b00111010111 : out <= 16'sb00000000_11111101; // 0.99210
        11'b00111011000 : out <= 16'sb00000000_11111110; // 0.99248
        11'b00111011001 : out <= 16'sb00000000_11111110; // 0.99285
        11'b00111011010 : out <= 16'sb00000000_11111110; // 0.99321
        11'b00111011011 : out <= 16'sb00000000_11111110; // 0.99356
        11'b00111011100 : out <= 16'sb00000000_11111110; // 0.99391
        11'b00111011101 : out <= 16'sb00000000_11111110; // 0.99424
        11'b00111011110 : out <= 16'sb00000000_11111110; // 0.99456
        11'b00111011111 : out <= 16'sb00000000_11111110; // 0.99488
        11'b00111100000 : out <= 16'sb00000000_11111110; // 0.99518
        11'b00111100001 : out <= 16'sb00000000_11111110; // 0.99548
        11'b00111100010 : out <= 16'sb00000000_11111110; // 0.99577
        11'b00111100011 : out <= 16'sb00000000_11111110; // 0.99604
        11'b00111100100 : out <= 16'sb00000000_11111111; // 0.99631
        11'b00111100101 : out <= 16'sb00000000_11111111; // 0.99657
        11'b00111100110 : out <= 16'sb00000000_11111111; // 0.99682
        11'b00111100111 : out <= 16'sb00000000_11111111; // 0.99706
        11'b00111101000 : out <= 16'sb00000000_11111111; // 0.99729
        11'b00111101001 : out <= 16'sb00000000_11111111; // 0.99751
        11'b00111101010 : out <= 16'sb00000000_11111111; // 0.99772
        11'b00111101011 : out <= 16'sb00000000_11111111; // 0.99793
        11'b00111101100 : out <= 16'sb00000000_11111111; // 0.99812
        11'b00111101101 : out <= 16'sb00000000_11111111; // 0.99830
        11'b00111101110 : out <= 16'sb00000000_11111111; // 0.99848
        11'b00111101111 : out <= 16'sb00000000_11111111; // 0.99864
        11'b00111110000 : out <= 16'sb00000000_11111111; // 0.99880
        11'b00111110001 : out <= 16'sb00000000_11111111; // 0.99894
        11'b00111110010 : out <= 16'sb00000000_11111111; // 0.99908
        11'b00111110011 : out <= 16'sb00000000_11111111; // 0.99920
        11'b00111110100 : out <= 16'sb00000000_11111111; // 0.99932
        11'b00111110101 : out <= 16'sb00000000_11111111; // 0.99943
        11'b00111110110 : out <= 16'sb00000000_11111111; // 0.99953
        11'b00111110111 : out <= 16'sb00000000_11111111; // 0.99962
        11'b00111111000 : out <= 16'sb00000000_11111111; // 0.99970
        11'b00111111001 : out <= 16'sb00000000_11111111; // 0.99977
        11'b00111111010 : out <= 16'sb00000000_11111111; // 0.99983
        11'b00111111011 : out <= 16'sb00000000_11111111; // 0.99988
        11'b00111111100 : out <= 16'sb00000000_11111111; // 0.99992
        11'b00111111101 : out <= 16'sb00000000_11111111; // 0.99996
        11'b00111111110 : out <= 16'sb00000000_11111111; // 0.99998
        11'b00111111111 : out <= 16'sb00000000_11111111; // 1.00000
        11'b01000000000 : out <= 16'sb00000001_00000000; // 1.00000
        11'b01000000001 : out <= 16'sb00000000_11111111; // 1.00000
        11'b01000000010 : out <= 16'sb00000000_11111111; // 0.99998
        11'b01000000011 : out <= 16'sb00000000_11111111; // 0.99996
        11'b01000000100 : out <= 16'sb00000000_11111111; // 0.99992
        11'b01000000101 : out <= 16'sb00000000_11111111; // 0.99988
        11'b01000000110 : out <= 16'sb00000000_11111111; // 0.99983
        11'b01000000111 : out <= 16'sb00000000_11111111; // 0.99977
        11'b01000001000 : out <= 16'sb00000000_11111111; // 0.99970
        11'b01000001001 : out <= 16'sb00000000_11111111; // 0.99962
        11'b01000001010 : out <= 16'sb00000000_11111111; // 0.99953
        11'b01000001011 : out <= 16'sb00000000_11111111; // 0.99943
        11'b01000001100 : out <= 16'sb00000000_11111111; // 0.99932
        11'b01000001101 : out <= 16'sb00000000_11111111; // 0.99920
        11'b01000001110 : out <= 16'sb00000000_11111111; // 0.99908
        11'b01000001111 : out <= 16'sb00000000_11111111; // 0.99894
        11'b01000010000 : out <= 16'sb00000000_11111111; // 0.99880
        11'b01000010001 : out <= 16'sb00000000_11111111; // 0.99864
        11'b01000010010 : out <= 16'sb00000000_11111111; // 0.99848
        11'b01000010011 : out <= 16'sb00000000_11111111; // 0.99830
        11'b01000010100 : out <= 16'sb00000000_11111111; // 0.99812
        11'b01000010101 : out <= 16'sb00000000_11111111; // 0.99793
        11'b01000010110 : out <= 16'sb00000000_11111111; // 0.99772
        11'b01000010111 : out <= 16'sb00000000_11111111; // 0.99751
        11'b01000011000 : out <= 16'sb00000000_11111111; // 0.99729
        11'b01000011001 : out <= 16'sb00000000_11111111; // 0.99706
        11'b01000011010 : out <= 16'sb00000000_11111111; // 0.99682
        11'b01000011011 : out <= 16'sb00000000_11111111; // 0.99657
        11'b01000011100 : out <= 16'sb00000000_11111111; // 0.99631
        11'b01000011101 : out <= 16'sb00000000_11111110; // 0.99604
        11'b01000011110 : out <= 16'sb00000000_11111110; // 0.99577
        11'b01000011111 : out <= 16'sb00000000_11111110; // 0.99548
        11'b01000100000 : out <= 16'sb00000000_11111110; // 0.99518
        11'b01000100001 : out <= 16'sb00000000_11111110; // 0.99488
        11'b01000100010 : out <= 16'sb00000000_11111110; // 0.99456
        11'b01000100011 : out <= 16'sb00000000_11111110; // 0.99424
        11'b01000100100 : out <= 16'sb00000000_11111110; // 0.99391
        11'b01000100101 : out <= 16'sb00000000_11111110; // 0.99356
        11'b01000100110 : out <= 16'sb00000000_11111110; // 0.99321
        11'b01000100111 : out <= 16'sb00000000_11111110; // 0.99285
        11'b01000101000 : out <= 16'sb00000000_11111110; // 0.99248
        11'b01000101001 : out <= 16'sb00000000_11111101; // 0.99210
        11'b01000101010 : out <= 16'sb00000000_11111101; // 0.99171
        11'b01000101011 : out <= 16'sb00000000_11111101; // 0.99131
        11'b01000101100 : out <= 16'sb00000000_11111101; // 0.99090
        11'b01000101101 : out <= 16'sb00000000_11111101; // 0.99049
        11'b01000101110 : out <= 16'sb00000000_11111101; // 0.99006
        11'b01000101111 : out <= 16'sb00000000_11111101; // 0.98962
        11'b01000110000 : out <= 16'sb00000000_11111101; // 0.98918
        11'b01000110001 : out <= 16'sb00000000_11111101; // 0.98872
        11'b01000110010 : out <= 16'sb00000000_11111100; // 0.98826
        11'b01000110011 : out <= 16'sb00000000_11111100; // 0.98778
        11'b01000110100 : out <= 16'sb00000000_11111100; // 0.98730
        11'b01000110101 : out <= 16'sb00000000_11111100; // 0.98681
        11'b01000110110 : out <= 16'sb00000000_11111100; // 0.98631
        11'b01000110111 : out <= 16'sb00000000_11111100; // 0.98580
        11'b01000111000 : out <= 16'sb00000000_11111100; // 0.98528
        11'b01000111001 : out <= 16'sb00000000_11111100; // 0.98475
        11'b01000111010 : out <= 16'sb00000000_11111011; // 0.98421
        11'b01000111011 : out <= 16'sb00000000_11111011; // 0.98366
        11'b01000111100 : out <= 16'sb00000000_11111011; // 0.98311
        11'b01000111101 : out <= 16'sb00000000_11111011; // 0.98254
        11'b01000111110 : out <= 16'sb00000000_11111011; // 0.98196
        11'b01000111111 : out <= 16'sb00000000_11111011; // 0.98138
        11'b01001000000 : out <= 16'sb00000000_11111011; // 0.98079
        11'b01001000001 : out <= 16'sb00000000_11111010; // 0.98018
        11'b01001000010 : out <= 16'sb00000000_11111010; // 0.97957
        11'b01001000011 : out <= 16'sb00000000_11111010; // 0.97895
        11'b01001000100 : out <= 16'sb00000000_11111010; // 0.97832
        11'b01001000101 : out <= 16'sb00000000_11111010; // 0.97768
        11'b01001000110 : out <= 16'sb00000000_11111010; // 0.97703
        11'b01001000111 : out <= 16'sb00000000_11111001; // 0.97637
        11'b01001001000 : out <= 16'sb00000000_11111001; // 0.97570
        11'b01001001001 : out <= 16'sb00000000_11111001; // 0.97503
        11'b01001001010 : out <= 16'sb00000000_11111001; // 0.97434
        11'b01001001011 : out <= 16'sb00000000_11111001; // 0.97364
        11'b01001001100 : out <= 16'sb00000000_11111001; // 0.97294
        11'b01001001101 : out <= 16'sb00000000_11111000; // 0.97223
        11'b01001001110 : out <= 16'sb00000000_11111000; // 0.97150
        11'b01001001111 : out <= 16'sb00000000_11111000; // 0.97077
        11'b01001010000 : out <= 16'sb00000000_11111000; // 0.97003
        11'b01001010001 : out <= 16'sb00000000_11111000; // 0.96928
        11'b01001010010 : out <= 16'sb00000000_11110111; // 0.96852
        11'b01001010011 : out <= 16'sb00000000_11110111; // 0.96775
        11'b01001010100 : out <= 16'sb00000000_11110111; // 0.96698
        11'b01001010101 : out <= 16'sb00000000_11110111; // 0.96619
        11'b01001010110 : out <= 16'sb00000000_11110111; // 0.96539
        11'b01001010111 : out <= 16'sb00000000_11110110; // 0.96459
        11'b01001011000 : out <= 16'sb00000000_11110110; // 0.96378
        11'b01001011001 : out <= 16'sb00000000_11110110; // 0.96295
        11'b01001011010 : out <= 16'sb00000000_11110110; // 0.96212
        11'b01001011011 : out <= 16'sb00000000_11110110; // 0.96128
        11'b01001011100 : out <= 16'sb00000000_11110101; // 0.96043
        11'b01001011101 : out <= 16'sb00000000_11110101; // 0.95957
        11'b01001011110 : out <= 16'sb00000000_11110101; // 0.95870
        11'b01001011111 : out <= 16'sb00000000_11110101; // 0.95783
        11'b01001100000 : out <= 16'sb00000000_11110100; // 0.95694
        11'b01001100001 : out <= 16'sb00000000_11110100; // 0.95605
        11'b01001100010 : out <= 16'sb00000000_11110100; // 0.95514
        11'b01001100011 : out <= 16'sb00000000_11110100; // 0.95423
        11'b01001100100 : out <= 16'sb00000000_11110100; // 0.95331
        11'b01001100101 : out <= 16'sb00000000_11110011; // 0.95238
        11'b01001100110 : out <= 16'sb00000000_11110011; // 0.95144
        11'b01001100111 : out <= 16'sb00000000_11110011; // 0.95049
        11'b01001101000 : out <= 16'sb00000000_11110011; // 0.94953
        11'b01001101001 : out <= 16'sb00000000_11110010; // 0.94856
        11'b01001101010 : out <= 16'sb00000000_11110010; // 0.94759
        11'b01001101011 : out <= 16'sb00000000_11110010; // 0.94660
        11'b01001101100 : out <= 16'sb00000000_11110010; // 0.94561
        11'b01001101101 : out <= 16'sb00000000_11110001; // 0.94460
        11'b01001101110 : out <= 16'sb00000000_11110001; // 0.94359
        11'b01001101111 : out <= 16'sb00000000_11110001; // 0.94257
        11'b01001110000 : out <= 16'sb00000000_11110001; // 0.94154
        11'b01001110001 : out <= 16'sb00000000_11110000; // 0.94051
        11'b01001110010 : out <= 16'sb00000000_11110000; // 0.93946
        11'b01001110011 : out <= 16'sb00000000_11110000; // 0.93840
        11'b01001110100 : out <= 16'sb00000000_11101111; // 0.93734
        11'b01001110101 : out <= 16'sb00000000_11101111; // 0.93627
        11'b01001110110 : out <= 16'sb00000000_11101111; // 0.93518
        11'b01001110111 : out <= 16'sb00000000_11101111; // 0.93409
        11'b01001111000 : out <= 16'sb00000000_11101110; // 0.93299
        11'b01001111001 : out <= 16'sb00000000_11101110; // 0.93188
        11'b01001111010 : out <= 16'sb00000000_11101110; // 0.93077
        11'b01001111011 : out <= 16'sb00000000_11101101; // 0.92964
        11'b01001111100 : out <= 16'sb00000000_11101101; // 0.92851
        11'b01001111101 : out <= 16'sb00000000_11101101; // 0.92736
        11'b01001111110 : out <= 16'sb00000000_11101101; // 0.92621
        11'b01001111111 : out <= 16'sb00000000_11101100; // 0.92505
        11'b01010000000 : out <= 16'sb00000000_11101100; // 0.92388
        11'b01010000001 : out <= 16'sb00000000_11101100; // 0.92270
        11'b01010000010 : out <= 16'sb00000000_11101011; // 0.92151
        11'b01010000011 : out <= 16'sb00000000_11101011; // 0.92032
        11'b01010000100 : out <= 16'sb00000000_11101011; // 0.91911
        11'b01010000101 : out <= 16'sb00000000_11101010; // 0.91790
        11'b01010000110 : out <= 16'sb00000000_11101010; // 0.91668
        11'b01010000111 : out <= 16'sb00000000_11101010; // 0.91545
        11'b01010001000 : out <= 16'sb00000000_11101010; // 0.91421
        11'b01010001001 : out <= 16'sb00000000_11101001; // 0.91296
        11'b01010001010 : out <= 16'sb00000000_11101001; // 0.91171
        11'b01010001011 : out <= 16'sb00000000_11101001; // 0.91044
        11'b01010001100 : out <= 16'sb00000000_11101000; // 0.90917
        11'b01010001101 : out <= 16'sb00000000_11101000; // 0.90789
        11'b01010001110 : out <= 16'sb00000000_11101000; // 0.90660
        11'b01010001111 : out <= 16'sb00000000_11100111; // 0.90530
        11'b01010010000 : out <= 16'sb00000000_11100111; // 0.90399
        11'b01010010001 : out <= 16'sb00000000_11100111; // 0.90267
        11'b01010010010 : out <= 16'sb00000000_11100110; // 0.90135
        11'b01010010011 : out <= 16'sb00000000_11100110; // 0.90002
        11'b01010010100 : out <= 16'sb00000000_11100110; // 0.89867
        11'b01010010101 : out <= 16'sb00000000_11100101; // 0.89732
        11'b01010010110 : out <= 16'sb00000000_11100101; // 0.89597
        11'b01010010111 : out <= 16'sb00000000_11100101; // 0.89460
        11'b01010011000 : out <= 16'sb00000000_11100100; // 0.89322
        11'b01010011001 : out <= 16'sb00000000_11100100; // 0.89184
        11'b01010011010 : out <= 16'sb00000000_11100011; // 0.89045
        11'b01010011011 : out <= 16'sb00000000_11100011; // 0.88905
        11'b01010011100 : out <= 16'sb00000000_11100011; // 0.88764
        11'b01010011101 : out <= 16'sb00000000_11100010; // 0.88622
        11'b01010011110 : out <= 16'sb00000000_11100010; // 0.88480
        11'b01010011111 : out <= 16'sb00000000_11100010; // 0.88336
        11'b01010100000 : out <= 16'sb00000000_11100001; // 0.88192
        11'b01010100001 : out <= 16'sb00000000_11100001; // 0.88047
        11'b01010100010 : out <= 16'sb00000000_11100001; // 0.87901
        11'b01010100011 : out <= 16'sb00000000_11100000; // 0.87755
        11'b01010100100 : out <= 16'sb00000000_11100000; // 0.87607
        11'b01010100101 : out <= 16'sb00000000_11011111; // 0.87459
        11'b01010100110 : out <= 16'sb00000000_11011111; // 0.87309
        11'b01010100111 : out <= 16'sb00000000_11011111; // 0.87160
        11'b01010101000 : out <= 16'sb00000000_11011110; // 0.87009
        11'b01010101001 : out <= 16'sb00000000_11011110; // 0.86857
        11'b01010101010 : out <= 16'sb00000000_11011101; // 0.86705
        11'b01010101011 : out <= 16'sb00000000_11011101; // 0.86551
        11'b01010101100 : out <= 16'sb00000000_11011101; // 0.86397
        11'b01010101101 : out <= 16'sb00000000_11011100; // 0.86242
        11'b01010101110 : out <= 16'sb00000000_11011100; // 0.86087
        11'b01010101111 : out <= 16'sb00000000_11011011; // 0.85930
        11'b01010110000 : out <= 16'sb00000000_11011011; // 0.85773
        11'b01010110001 : out <= 16'sb00000000_11011011; // 0.85615
        11'b01010110010 : out <= 16'sb00000000_11011010; // 0.85456
        11'b01010110011 : out <= 16'sb00000000_11011010; // 0.85296
        11'b01010110100 : out <= 16'sb00000000_11011001; // 0.85136
        11'b01010110101 : out <= 16'sb00000000_11011001; // 0.84974
        11'b01010110110 : out <= 16'sb00000000_11011001; // 0.84812
        11'b01010110111 : out <= 16'sb00000000_11011000; // 0.84649
        11'b01010111000 : out <= 16'sb00000000_11011000; // 0.84485
        11'b01010111001 : out <= 16'sb00000000_11010111; // 0.84321
        11'b01010111010 : out <= 16'sb00000000_11010111; // 0.84155
        11'b01010111011 : out <= 16'sb00000000_11010111; // 0.83989
        11'b01010111100 : out <= 16'sb00000000_11010110; // 0.83822
        11'b01010111101 : out <= 16'sb00000000_11010110; // 0.83655
        11'b01010111110 : out <= 16'sb00000000_11010101; // 0.83486
        11'b01010111111 : out <= 16'sb00000000_11010101; // 0.83317
        11'b01011000000 : out <= 16'sb00000000_11010100; // 0.83147
        11'b01011000001 : out <= 16'sb00000000_11010100; // 0.82976
        11'b01011000010 : out <= 16'sb00000000_11010011; // 0.82805
        11'b01011000011 : out <= 16'sb00000000_11010011; // 0.82632
        11'b01011000100 : out <= 16'sb00000000_11010011; // 0.82459
        11'b01011000101 : out <= 16'sb00000000_11010010; // 0.82285
        11'b01011000110 : out <= 16'sb00000000_11010010; // 0.82110
        11'b01011000111 : out <= 16'sb00000000_11010001; // 0.81935
        11'b01011001000 : out <= 16'sb00000000_11010001; // 0.81758
        11'b01011001001 : out <= 16'sb00000000_11010000; // 0.81581
        11'b01011001010 : out <= 16'sb00000000_11010000; // 0.81404
        11'b01011001011 : out <= 16'sb00000000_11001111; // 0.81225
        11'b01011001100 : out <= 16'sb00000000_11001111; // 0.81046
        11'b01011001101 : out <= 16'sb00000000_11001111; // 0.80866
        11'b01011001110 : out <= 16'sb00000000_11001110; // 0.80685
        11'b01011001111 : out <= 16'sb00000000_11001110; // 0.80503
        11'b01011010000 : out <= 16'sb00000000_11001101; // 0.80321
        11'b01011010001 : out <= 16'sb00000000_11001101; // 0.80138
        11'b01011010010 : out <= 16'sb00000000_11001100; // 0.79954
        11'b01011010011 : out <= 16'sb00000000_11001100; // 0.79769
        11'b01011010100 : out <= 16'sb00000000_11001011; // 0.79584
        11'b01011010101 : out <= 16'sb00000000_11001011; // 0.79398
        11'b01011010110 : out <= 16'sb00000000_11001010; // 0.79211
        11'b01011010111 : out <= 16'sb00000000_11001010; // 0.79023
        11'b01011011000 : out <= 16'sb00000000_11001001; // 0.78835
        11'b01011011001 : out <= 16'sb00000000_11001001; // 0.78646
        11'b01011011010 : out <= 16'sb00000000_11001000; // 0.78456
        11'b01011011011 : out <= 16'sb00000000_11001000; // 0.78265
        11'b01011011100 : out <= 16'sb00000000_11000111; // 0.78074
        11'b01011011101 : out <= 16'sb00000000_11000111; // 0.77882
        11'b01011011110 : out <= 16'sb00000000_11000110; // 0.77689
        11'b01011011111 : out <= 16'sb00000000_11000110; // 0.77495
        11'b01011100000 : out <= 16'sb00000000_11000101; // 0.77301
        11'b01011100001 : out <= 16'sb00000000_11000101; // 0.77106
        11'b01011100010 : out <= 16'sb00000000_11000100; // 0.76910
        11'b01011100011 : out <= 16'sb00000000_11000100; // 0.76714
        11'b01011100100 : out <= 16'sb00000000_11000011; // 0.76517
        11'b01011100101 : out <= 16'sb00000000_11000011; // 0.76319
        11'b01011100110 : out <= 16'sb00000000_11000010; // 0.76120
        11'b01011100111 : out <= 16'sb00000000_11000010; // 0.75921
        11'b01011101000 : out <= 16'sb00000000_11000001; // 0.75721
        11'b01011101001 : out <= 16'sb00000000_11000001; // 0.75520
        11'b01011101010 : out <= 16'sb00000000_11000000; // 0.75319
        11'b01011101011 : out <= 16'sb00000000_11000000; // 0.75117
        11'b01011101100 : out <= 16'sb00000000_10111111; // 0.74914
        11'b01011101101 : out <= 16'sb00000000_10111111; // 0.74710
        11'b01011101110 : out <= 16'sb00000000_10111110; // 0.74506
        11'b01011101111 : out <= 16'sb00000000_10111110; // 0.74301
        11'b01011110000 : out <= 16'sb00000000_10111101; // 0.74095
        11'b01011110001 : out <= 16'sb00000000_10111101; // 0.73889
        11'b01011110010 : out <= 16'sb00000000_10111100; // 0.73682
        11'b01011110011 : out <= 16'sb00000000_10111100; // 0.73474
        11'b01011110100 : out <= 16'sb00000000_10111011; // 0.73265
        11'b01011110101 : out <= 16'sb00000000_10111011; // 0.73056
        11'b01011110110 : out <= 16'sb00000000_10111010; // 0.72846
        11'b01011110111 : out <= 16'sb00000000_10111001; // 0.72636
        11'b01011111000 : out <= 16'sb00000000_10111001; // 0.72425
        11'b01011111001 : out <= 16'sb00000000_10111000; // 0.72213
        11'b01011111010 : out <= 16'sb00000000_10111000; // 0.72000
        11'b01011111011 : out <= 16'sb00000000_10110111; // 0.71787
        11'b01011111100 : out <= 16'sb00000000_10110111; // 0.71573
        11'b01011111101 : out <= 16'sb00000000_10110110; // 0.71358
        11'b01011111110 : out <= 16'sb00000000_10110110; // 0.71143
        11'b01011111111 : out <= 16'sb00000000_10110101; // 0.70927
        11'b01100000000 : out <= 16'sb00000000_10110101; // 0.70711
        11'b01100000001 : out <= 16'sb00000000_10110100; // 0.70493
        11'b01100000010 : out <= 16'sb00000000_10110011; // 0.70275
        11'b01100000011 : out <= 16'sb00000000_10110011; // 0.70057
        11'b01100000100 : out <= 16'sb00000000_10110010; // 0.69838
        11'b01100000101 : out <= 16'sb00000000_10110010; // 0.69618
        11'b01100000110 : out <= 16'sb00000000_10110001; // 0.69397
        11'b01100000111 : out <= 16'sb00000000_10110001; // 0.69176
        11'b01100001000 : out <= 16'sb00000000_10110000; // 0.68954
        11'b01100001001 : out <= 16'sb00000000_10101111; // 0.68732
        11'b01100001010 : out <= 16'sb00000000_10101111; // 0.68508
        11'b01100001011 : out <= 16'sb00000000_10101110; // 0.68285
        11'b01100001100 : out <= 16'sb00000000_10101110; // 0.68060
        11'b01100001101 : out <= 16'sb00000000_10101101; // 0.67835
        11'b01100001110 : out <= 16'sb00000000_10101101; // 0.67609
        11'b01100001111 : out <= 16'sb00000000_10101100; // 0.67383
        11'b01100010000 : out <= 16'sb00000000_10101011; // 0.67156
        11'b01100010001 : out <= 16'sb00000000_10101011; // 0.66928
        11'b01100010010 : out <= 16'sb00000000_10101010; // 0.66700
        11'b01100010011 : out <= 16'sb00000000_10101010; // 0.66471
        11'b01100010100 : out <= 16'sb00000000_10101001; // 0.66242
        11'b01100010101 : out <= 16'sb00000000_10101000; // 0.66011
        11'b01100010110 : out <= 16'sb00000000_10101000; // 0.65781
        11'b01100010111 : out <= 16'sb00000000_10100111; // 0.65549
        11'b01100011000 : out <= 16'sb00000000_10100111; // 0.65317
        11'b01100011001 : out <= 16'sb00000000_10100110; // 0.65085
        11'b01100011010 : out <= 16'sb00000000_10100110; // 0.64851
        11'b01100011011 : out <= 16'sb00000000_10100101; // 0.64618
        11'b01100011100 : out <= 16'sb00000000_10100100; // 0.64383
        11'b01100011101 : out <= 16'sb00000000_10100100; // 0.64148
        11'b01100011110 : out <= 16'sb00000000_10100011; // 0.63912
        11'b01100011111 : out <= 16'sb00000000_10100011; // 0.63676
        11'b01100100000 : out <= 16'sb00000000_10100010; // 0.63439
        11'b01100100001 : out <= 16'sb00000000_10100001; // 0.63202
        11'b01100100010 : out <= 16'sb00000000_10100001; // 0.62964
        11'b01100100011 : out <= 16'sb00000000_10100000; // 0.62725
        11'b01100100100 : out <= 16'sb00000000_10011111; // 0.62486
        11'b01100100101 : out <= 16'sb00000000_10011111; // 0.62246
        11'b01100100110 : out <= 16'sb00000000_10011110; // 0.62006
        11'b01100100111 : out <= 16'sb00000000_10011110; // 0.61765
        11'b01100101000 : out <= 16'sb00000000_10011101; // 0.61523
        11'b01100101001 : out <= 16'sb00000000_10011100; // 0.61281
        11'b01100101010 : out <= 16'sb00000000_10011100; // 0.61038
        11'b01100101011 : out <= 16'sb00000000_10011011; // 0.60795
        11'b01100101100 : out <= 16'sb00000000_10011011; // 0.60551
        11'b01100101101 : out <= 16'sb00000000_10011010; // 0.60307
        11'b01100101110 : out <= 16'sb00000000_10011001; // 0.60062
        11'b01100101111 : out <= 16'sb00000000_10011001; // 0.59816
        11'b01100110000 : out <= 16'sb00000000_10011000; // 0.59570
        11'b01100110001 : out <= 16'sb00000000_10010111; // 0.59323
        11'b01100110010 : out <= 16'sb00000000_10010111; // 0.59076
        11'b01100110011 : out <= 16'sb00000000_10010110; // 0.58828
        11'b01100110100 : out <= 16'sb00000000_10010101; // 0.58580
        11'b01100110101 : out <= 16'sb00000000_10010101; // 0.58331
        11'b01100110110 : out <= 16'sb00000000_10010100; // 0.58081
        11'b01100110111 : out <= 16'sb00000000_10010100; // 0.57831
        11'b01100111000 : out <= 16'sb00000000_10010011; // 0.57581
        11'b01100111001 : out <= 16'sb00000000_10010010; // 0.57330
        11'b01100111010 : out <= 16'sb00000000_10010010; // 0.57078
        11'b01100111011 : out <= 16'sb00000000_10010001; // 0.56826
        11'b01100111100 : out <= 16'sb00000000_10010000; // 0.56573
        11'b01100111101 : out <= 16'sb00000000_10010000; // 0.56320
        11'b01100111110 : out <= 16'sb00000000_10001111; // 0.56066
        11'b01100111111 : out <= 16'sb00000000_10001110; // 0.55812
        11'b01101000000 : out <= 16'sb00000000_10001110; // 0.55557
        11'b01101000001 : out <= 16'sb00000000_10001101; // 0.55302
        11'b01101000010 : out <= 16'sb00000000_10001100; // 0.55046
        11'b01101000011 : out <= 16'sb00000000_10001100; // 0.54789
        11'b01101000100 : out <= 16'sb00000000_10001011; // 0.54532
        11'b01101000101 : out <= 16'sb00000000_10001010; // 0.54275
        11'b01101000110 : out <= 16'sb00000000_10001010; // 0.54017
        11'b01101000111 : out <= 16'sb00000000_10001001; // 0.53759
        11'b01101001000 : out <= 16'sb00000000_10001000; // 0.53500
        11'b01101001001 : out <= 16'sb00000000_10001000; // 0.53240
        11'b01101001010 : out <= 16'sb00000000_10000111; // 0.52980
        11'b01101001011 : out <= 16'sb00000000_10000110; // 0.52720
        11'b01101001100 : out <= 16'sb00000000_10000110; // 0.52459
        11'b01101001101 : out <= 16'sb00000000_10000101; // 0.52198
        11'b01101001110 : out <= 16'sb00000000_10000100; // 0.51936
        11'b01101001111 : out <= 16'sb00000000_10000100; // 0.51673
        11'b01101010000 : out <= 16'sb00000000_10000011; // 0.51410
        11'b01101010001 : out <= 16'sb00000000_10000010; // 0.51147
        11'b01101010010 : out <= 16'sb00000000_10000010; // 0.50883
        11'b01101010011 : out <= 16'sb00000000_10000001; // 0.50619
        11'b01101010100 : out <= 16'sb00000000_10000000; // 0.50354
        11'b01101010101 : out <= 16'sb00000000_10000000; // 0.50089
        11'b01101010110 : out <= 16'sb00000000_01111111; // 0.49823
        11'b01101010111 : out <= 16'sb00000000_01111110; // 0.49557
        11'b01101011000 : out <= 16'sb00000000_01111110; // 0.49290
        11'b01101011001 : out <= 16'sb00000000_01111101; // 0.49023
        11'b01101011010 : out <= 16'sb00000000_01111100; // 0.48755
        11'b01101011011 : out <= 16'sb00000000_01111100; // 0.48487
        11'b01101011100 : out <= 16'sb00000000_01111011; // 0.48218
        11'b01101011101 : out <= 16'sb00000000_01111010; // 0.47949
        11'b01101011110 : out <= 16'sb00000000_01111010; // 0.47680
        11'b01101011111 : out <= 16'sb00000000_01111001; // 0.47410
        11'b01101100000 : out <= 16'sb00000000_01111000; // 0.47140
        11'b01101100001 : out <= 16'sb00000000_01110111; // 0.46869
        11'b01101100010 : out <= 16'sb00000000_01110111; // 0.46598
        11'b01101100011 : out <= 16'sb00000000_01110110; // 0.46326
        11'b01101100100 : out <= 16'sb00000000_01110101; // 0.46054
        11'b01101100101 : out <= 16'sb00000000_01110101; // 0.45781
        11'b01101100110 : out <= 16'sb00000000_01110100; // 0.45508
        11'b01101100111 : out <= 16'sb00000000_01110011; // 0.45235
        11'b01101101000 : out <= 16'sb00000000_01110011; // 0.44961
        11'b01101101001 : out <= 16'sb00000000_01110010; // 0.44687
        11'b01101101010 : out <= 16'sb00000000_01110001; // 0.44412
        11'b01101101011 : out <= 16'sb00000000_01110000; // 0.44137
        11'b01101101100 : out <= 16'sb00000000_01110000; // 0.43862
        11'b01101101101 : out <= 16'sb00000000_01101111; // 0.43586
        11'b01101101110 : out <= 16'sb00000000_01101110; // 0.43309
        11'b01101101111 : out <= 16'sb00000000_01101110; // 0.43033
        11'b01101110000 : out <= 16'sb00000000_01101101; // 0.42756
        11'b01101110001 : out <= 16'sb00000000_01101100; // 0.42478
        11'b01101110010 : out <= 16'sb00000000_01101100; // 0.42200
        11'b01101110011 : out <= 16'sb00000000_01101011; // 0.41922
        11'b01101110100 : out <= 16'sb00000000_01101010; // 0.41643
        11'b01101110101 : out <= 16'sb00000000_01101001; // 0.41364
        11'b01101110110 : out <= 16'sb00000000_01101001; // 0.41084
        11'b01101110111 : out <= 16'sb00000000_01101000; // 0.40804
        11'b01101111000 : out <= 16'sb00000000_01100111; // 0.40524
        11'b01101111001 : out <= 16'sb00000000_01100111; // 0.40243
        11'b01101111010 : out <= 16'sb00000000_01100110; // 0.39962
        11'b01101111011 : out <= 16'sb00000000_01100101; // 0.39681
        11'b01101111100 : out <= 16'sb00000000_01100100; // 0.39399
        11'b01101111101 : out <= 16'sb00000000_01100100; // 0.39117
        11'b01101111110 : out <= 16'sb00000000_01100011; // 0.38835
        11'b01101111111 : out <= 16'sb00000000_01100010; // 0.38552
        11'b01110000000 : out <= 16'sb00000000_01100001; // 0.38268
        11'b01110000001 : out <= 16'sb00000000_01100001; // 0.37985
        11'b01110000010 : out <= 16'sb00000000_01100000; // 0.37701
        11'b01110000011 : out <= 16'sb00000000_01011111; // 0.37416
        11'b01110000100 : out <= 16'sb00000000_01011111; // 0.37132
        11'b01110000101 : out <= 16'sb00000000_01011110; // 0.36847
        11'b01110000110 : out <= 16'sb00000000_01011101; // 0.36561
        11'b01110000111 : out <= 16'sb00000000_01011100; // 0.36276
        11'b01110001000 : out <= 16'sb00000000_01011100; // 0.35990
        11'b01110001001 : out <= 16'sb00000000_01011011; // 0.35703
        11'b01110001010 : out <= 16'sb00000000_01011010; // 0.35416
        11'b01110001011 : out <= 16'sb00000000_01011001; // 0.35129
        11'b01110001100 : out <= 16'sb00000000_01011001; // 0.34842
        11'b01110001101 : out <= 16'sb00000000_01011000; // 0.34554
        11'b01110001110 : out <= 16'sb00000000_01010111; // 0.34266
        11'b01110001111 : out <= 16'sb00000000_01010110; // 0.33978
        11'b01110010000 : out <= 16'sb00000000_01010110; // 0.33689
        11'b01110010001 : out <= 16'sb00000000_01010101; // 0.33400
        11'b01110010010 : out <= 16'sb00000000_01010100; // 0.33111
        11'b01110010011 : out <= 16'sb00000000_01010100; // 0.32821
        11'b01110010100 : out <= 16'sb00000000_01010011; // 0.32531
        11'b01110010101 : out <= 16'sb00000000_01010010; // 0.32241
        11'b01110010110 : out <= 16'sb00000000_01010001; // 0.31950
        11'b01110010111 : out <= 16'sb00000000_01010001; // 0.31659
        11'b01110011000 : out <= 16'sb00000000_01010000; // 0.31368
        11'b01110011001 : out <= 16'sb00000000_01001111; // 0.31077
        11'b01110011010 : out <= 16'sb00000000_01001110; // 0.30785
        11'b01110011011 : out <= 16'sb00000000_01001110; // 0.30493
        11'b01110011100 : out <= 16'sb00000000_01001101; // 0.30201
        11'b01110011101 : out <= 16'sb00000000_01001100; // 0.29908
        11'b01110011110 : out <= 16'sb00000000_01001011; // 0.29615
        11'b01110011111 : out <= 16'sb00000000_01001011; // 0.29322
        11'b01110100000 : out <= 16'sb00000000_01001010; // 0.29028
        11'b01110100001 : out <= 16'sb00000000_01001001; // 0.28735
        11'b01110100010 : out <= 16'sb00000000_01001000; // 0.28441
        11'b01110100011 : out <= 16'sb00000000_01001000; // 0.28146
        11'b01110100100 : out <= 16'sb00000000_01000111; // 0.27852
        11'b01110100101 : out <= 16'sb00000000_01000110; // 0.27557
        11'b01110100110 : out <= 16'sb00000000_01000101; // 0.27262
        11'b01110100111 : out <= 16'sb00000000_01000101; // 0.26967
        11'b01110101000 : out <= 16'sb00000000_01000100; // 0.26671
        11'b01110101001 : out <= 16'sb00000000_01000011; // 0.26375
        11'b01110101010 : out <= 16'sb00000000_01000010; // 0.26079
        11'b01110101011 : out <= 16'sb00000000_01000010; // 0.25783
        11'b01110101100 : out <= 16'sb00000000_01000001; // 0.25487
        11'b01110101101 : out <= 16'sb00000000_01000000; // 0.25190
        11'b01110101110 : out <= 16'sb00000000_00111111; // 0.24893
        11'b01110101111 : out <= 16'sb00000000_00111110; // 0.24596
        11'b01110110000 : out <= 16'sb00000000_00111110; // 0.24298
        11'b01110110001 : out <= 16'sb00000000_00111101; // 0.24000
        11'b01110110010 : out <= 16'sb00000000_00111100; // 0.23702
        11'b01110110011 : out <= 16'sb00000000_00111011; // 0.23404
        11'b01110110100 : out <= 16'sb00000000_00111011; // 0.23106
        11'b01110110101 : out <= 16'sb00000000_00111010; // 0.22807
        11'b01110110110 : out <= 16'sb00000000_00111001; // 0.22508
        11'b01110110111 : out <= 16'sb00000000_00111000; // 0.22209
        11'b01110111000 : out <= 16'sb00000000_00111000; // 0.21910
        11'b01110111001 : out <= 16'sb00000000_00110111; // 0.21611
        11'b01110111010 : out <= 16'sb00000000_00110110; // 0.21311
        11'b01110111011 : out <= 16'sb00000000_00110101; // 0.21011
        11'b01110111100 : out <= 16'sb00000000_00110101; // 0.20711
        11'b01110111101 : out <= 16'sb00000000_00110100; // 0.20411
        11'b01110111110 : out <= 16'sb00000000_00110011; // 0.20110
        11'b01110111111 : out <= 16'sb00000000_00110010; // 0.19810
        11'b01111000000 : out <= 16'sb00000000_00110001; // 0.19509
        11'b01111000001 : out <= 16'sb00000000_00110001; // 0.19208
        11'b01111000010 : out <= 16'sb00000000_00110000; // 0.18907
        11'b01111000011 : out <= 16'sb00000000_00101111; // 0.18606
        11'b01111000100 : out <= 16'sb00000000_00101110; // 0.18304
        11'b01111000101 : out <= 16'sb00000000_00101110; // 0.18002
        11'b01111000110 : out <= 16'sb00000000_00101101; // 0.17700
        11'b01111000111 : out <= 16'sb00000000_00101100; // 0.17398
        11'b01111001000 : out <= 16'sb00000000_00101011; // 0.17096
        11'b01111001001 : out <= 16'sb00000000_00101010; // 0.16794
        11'b01111001010 : out <= 16'sb00000000_00101010; // 0.16491
        11'b01111001011 : out <= 16'sb00000000_00101001; // 0.16189
        11'b01111001100 : out <= 16'sb00000000_00101000; // 0.15886
        11'b01111001101 : out <= 16'sb00000000_00100111; // 0.15583
        11'b01111001110 : out <= 16'sb00000000_00100111; // 0.15280
        11'b01111001111 : out <= 16'sb00000000_00100110; // 0.14976
        11'b01111010000 : out <= 16'sb00000000_00100101; // 0.14673
        11'b01111010001 : out <= 16'sb00000000_00100100; // 0.14370
        11'b01111010010 : out <= 16'sb00000000_00100100; // 0.14066
        11'b01111010011 : out <= 16'sb00000000_00100011; // 0.13762
        11'b01111010100 : out <= 16'sb00000000_00100010; // 0.13458
        11'b01111010101 : out <= 16'sb00000000_00100001; // 0.13154
        11'b01111010110 : out <= 16'sb00000000_00100000; // 0.12850
        11'b01111010111 : out <= 16'sb00000000_00100000; // 0.12545
        11'b01111011000 : out <= 16'sb00000000_00011111; // 0.12241
        11'b01111011001 : out <= 16'sb00000000_00011110; // 0.11937
        11'b01111011010 : out <= 16'sb00000000_00011101; // 0.11632
        11'b01111011011 : out <= 16'sb00000000_00011100; // 0.11327
        11'b01111011100 : out <= 16'sb00000000_00011100; // 0.11022
        11'b01111011101 : out <= 16'sb00000000_00011011; // 0.10717
        11'b01111011110 : out <= 16'sb00000000_00011010; // 0.10412
        11'b01111011111 : out <= 16'sb00000000_00011001; // 0.10107
        11'b01111100000 : out <= 16'sb00000000_00011001; // 0.09802
        11'b01111100001 : out <= 16'sb00000000_00011000; // 0.09496
        11'b01111100010 : out <= 16'sb00000000_00010111; // 0.09191
        11'b01111100011 : out <= 16'sb00000000_00010110; // 0.08885
        11'b01111100100 : out <= 16'sb00000000_00010101; // 0.08580
        11'b01111100101 : out <= 16'sb00000000_00010101; // 0.08274
        11'b01111100110 : out <= 16'sb00000000_00010100; // 0.07968
        11'b01111100111 : out <= 16'sb00000000_00010011; // 0.07662
        11'b01111101000 : out <= 16'sb00000000_00010010; // 0.07356
        11'b01111101001 : out <= 16'sb00000000_00010010; // 0.07050
        11'b01111101010 : out <= 16'sb00000000_00010001; // 0.06744
        11'b01111101011 : out <= 16'sb00000000_00010000; // 0.06438
        11'b01111101100 : out <= 16'sb00000000_00001111; // 0.06132
        11'b01111101101 : out <= 16'sb00000000_00001110; // 0.05826
        11'b01111101110 : out <= 16'sb00000000_00001110; // 0.05520
        11'b01111101111 : out <= 16'sb00000000_00001101; // 0.05213
        11'b01111110000 : out <= 16'sb00000000_00001100; // 0.04907
        11'b01111110001 : out <= 16'sb00000000_00001011; // 0.04600
        11'b01111110010 : out <= 16'sb00000000_00001010; // 0.04294
        11'b01111110011 : out <= 16'sb00000000_00001010; // 0.03987
        11'b01111110100 : out <= 16'sb00000000_00001001; // 0.03681
        11'b01111110101 : out <= 16'sb00000000_00001000; // 0.03374
        11'b01111110110 : out <= 16'sb00000000_00000111; // 0.03067
        11'b01111110111 : out <= 16'sb00000000_00000111; // 0.02761
        11'b01111111000 : out <= 16'sb00000000_00000110; // 0.02454
        11'b01111111001 : out <= 16'sb00000000_00000101; // 0.02147
        11'b01111111010 : out <= 16'sb00000000_00000100; // 0.01841
        11'b01111111011 : out <= 16'sb00000000_00000011; // 0.01534
        11'b01111111100 : out <= 16'sb00000000_00000011; // 0.01227
        11'b01111111101 : out <= 16'sb00000000_00000010; // 0.00920
        11'b01111111110 : out <= 16'sb00000000_00000001; // 0.00614
        11'b01111111111 : out <= 16'sb00000000_00000000; // 0.00307
        11'b10000000000 : out <= 16'sb00000000_00000000; // 0.00000
        11'b10000000001 : out <= 16'sb00000000_00000000; // -0.00307
        11'b10000000010 : out <= 16'sb11111111_11111111; // -0.00614
        11'b10000000011 : out <= 16'sb11111111_11111110; // -0.00920
        11'b10000000100 : out <= 16'sb11111111_11111101; // -0.01227
        11'b10000000101 : out <= 16'sb11111111_11111101; // -0.01534
        11'b10000000110 : out <= 16'sb11111111_11111100; // -0.01841
        11'b10000000111 : out <= 16'sb11111111_11111011; // -0.02147
        11'b10000001000 : out <= 16'sb11111111_11111010; // -0.02454
        11'b10000001001 : out <= 16'sb11111111_11111001; // -0.02761
        11'b10000001010 : out <= 16'sb11111111_11111001; // -0.03067
        11'b10000001011 : out <= 16'sb11111111_11111000; // -0.03374
        11'b10000001100 : out <= 16'sb11111111_11110111; // -0.03681
        11'b10000001101 : out <= 16'sb11111111_11110110; // -0.03987
        11'b10000001110 : out <= 16'sb11111111_11110110; // -0.04294
        11'b10000001111 : out <= 16'sb11111111_11110101; // -0.04600
        11'b10000010000 : out <= 16'sb11111111_11110100; // -0.04907
        11'b10000010001 : out <= 16'sb11111111_11110011; // -0.05213
        11'b10000010010 : out <= 16'sb11111111_11110010; // -0.05520
        11'b10000010011 : out <= 16'sb11111111_11110010; // -0.05826
        11'b10000010100 : out <= 16'sb11111111_11110001; // -0.06132
        11'b10000010101 : out <= 16'sb11111111_11110000; // -0.06438
        11'b10000010110 : out <= 16'sb11111111_11101111; // -0.06744
        11'b10000010111 : out <= 16'sb11111111_11101110; // -0.07050
        11'b10000011000 : out <= 16'sb11111111_11101110; // -0.07356
        11'b10000011001 : out <= 16'sb11111111_11101101; // -0.07662
        11'b10000011010 : out <= 16'sb11111111_11101100; // -0.07968
        11'b10000011011 : out <= 16'sb11111111_11101011; // -0.08274
        11'b10000011100 : out <= 16'sb11111111_11101011; // -0.08580
        11'b10000011101 : out <= 16'sb11111111_11101010; // -0.08885
        11'b10000011110 : out <= 16'sb11111111_11101001; // -0.09191
        11'b10000011111 : out <= 16'sb11111111_11101000; // -0.09496
        11'b10000100000 : out <= 16'sb11111111_11100111; // -0.09802
        11'b10000100001 : out <= 16'sb11111111_11100111; // -0.10107
        11'b10000100010 : out <= 16'sb11111111_11100110; // -0.10412
        11'b10000100011 : out <= 16'sb11111111_11100101; // -0.10717
        11'b10000100100 : out <= 16'sb11111111_11100100; // -0.11022
        11'b10000100101 : out <= 16'sb11111111_11100100; // -0.11327
        11'b10000100110 : out <= 16'sb11111111_11100011; // -0.11632
        11'b10000100111 : out <= 16'sb11111111_11100010; // -0.11937
        11'b10000101000 : out <= 16'sb11111111_11100001; // -0.12241
        11'b10000101001 : out <= 16'sb11111111_11100000; // -0.12545
        11'b10000101010 : out <= 16'sb11111111_11100000; // -0.12850
        11'b10000101011 : out <= 16'sb11111111_11011111; // -0.13154
        11'b10000101100 : out <= 16'sb11111111_11011110; // -0.13458
        11'b10000101101 : out <= 16'sb11111111_11011101; // -0.13762
        11'b10000101110 : out <= 16'sb11111111_11011100; // -0.14066
        11'b10000101111 : out <= 16'sb11111111_11011100; // -0.14370
        11'b10000110000 : out <= 16'sb11111111_11011011; // -0.14673
        11'b10000110001 : out <= 16'sb11111111_11011010; // -0.14976
        11'b10000110010 : out <= 16'sb11111111_11011001; // -0.15280
        11'b10000110011 : out <= 16'sb11111111_11011001; // -0.15583
        11'b10000110100 : out <= 16'sb11111111_11011000; // -0.15886
        11'b10000110101 : out <= 16'sb11111111_11010111; // -0.16189
        11'b10000110110 : out <= 16'sb11111111_11010110; // -0.16491
        11'b10000110111 : out <= 16'sb11111111_11010110; // -0.16794
        11'b10000111000 : out <= 16'sb11111111_11010101; // -0.17096
        11'b10000111001 : out <= 16'sb11111111_11010100; // -0.17398
        11'b10000111010 : out <= 16'sb11111111_11010011; // -0.17700
        11'b10000111011 : out <= 16'sb11111111_11010010; // -0.18002
        11'b10000111100 : out <= 16'sb11111111_11010010; // -0.18304
        11'b10000111101 : out <= 16'sb11111111_11010001; // -0.18606
        11'b10000111110 : out <= 16'sb11111111_11010000; // -0.18907
        11'b10000111111 : out <= 16'sb11111111_11001111; // -0.19208
        11'b10001000000 : out <= 16'sb11111111_11001111; // -0.19509
        11'b10001000001 : out <= 16'sb11111111_11001110; // -0.19810
        11'b10001000010 : out <= 16'sb11111111_11001101; // -0.20110
        11'b10001000011 : out <= 16'sb11111111_11001100; // -0.20411
        11'b10001000100 : out <= 16'sb11111111_11001011; // -0.20711
        11'b10001000101 : out <= 16'sb11111111_11001011; // -0.21011
        11'b10001000110 : out <= 16'sb11111111_11001010; // -0.21311
        11'b10001000111 : out <= 16'sb11111111_11001001; // -0.21611
        11'b10001001000 : out <= 16'sb11111111_11001000; // -0.21910
        11'b10001001001 : out <= 16'sb11111111_11001000; // -0.22209
        11'b10001001010 : out <= 16'sb11111111_11000111; // -0.22508
        11'b10001001011 : out <= 16'sb11111111_11000110; // -0.22807
        11'b10001001100 : out <= 16'sb11111111_11000101; // -0.23106
        11'b10001001101 : out <= 16'sb11111111_11000101; // -0.23404
        11'b10001001110 : out <= 16'sb11111111_11000100; // -0.23702
        11'b10001001111 : out <= 16'sb11111111_11000011; // -0.24000
        11'b10001010000 : out <= 16'sb11111111_11000010; // -0.24298
        11'b10001010001 : out <= 16'sb11111111_11000010; // -0.24596
        11'b10001010010 : out <= 16'sb11111111_11000001; // -0.24893
        11'b10001010011 : out <= 16'sb11111111_11000000; // -0.25190
        11'b10001010100 : out <= 16'sb11111111_10111111; // -0.25487
        11'b10001010101 : out <= 16'sb11111111_10111110; // -0.25783
        11'b10001010110 : out <= 16'sb11111111_10111110; // -0.26079
        11'b10001010111 : out <= 16'sb11111111_10111101; // -0.26375
        11'b10001011000 : out <= 16'sb11111111_10111100; // -0.26671
        11'b10001011001 : out <= 16'sb11111111_10111011; // -0.26967
        11'b10001011010 : out <= 16'sb11111111_10111011; // -0.27262
        11'b10001011011 : out <= 16'sb11111111_10111010; // -0.27557
        11'b10001011100 : out <= 16'sb11111111_10111001; // -0.27852
        11'b10001011101 : out <= 16'sb11111111_10111000; // -0.28146
        11'b10001011110 : out <= 16'sb11111111_10111000; // -0.28441
        11'b10001011111 : out <= 16'sb11111111_10110111; // -0.28735
        11'b10001100000 : out <= 16'sb11111111_10110110; // -0.29028
        11'b10001100001 : out <= 16'sb11111111_10110101; // -0.29322
        11'b10001100010 : out <= 16'sb11111111_10110101; // -0.29615
        11'b10001100011 : out <= 16'sb11111111_10110100; // -0.29908
        11'b10001100100 : out <= 16'sb11111111_10110011; // -0.30201
        11'b10001100101 : out <= 16'sb11111111_10110010; // -0.30493
        11'b10001100110 : out <= 16'sb11111111_10110010; // -0.30785
        11'b10001100111 : out <= 16'sb11111111_10110001; // -0.31077
        11'b10001101000 : out <= 16'sb11111111_10110000; // -0.31368
        11'b10001101001 : out <= 16'sb11111111_10101111; // -0.31659
        11'b10001101010 : out <= 16'sb11111111_10101111; // -0.31950
        11'b10001101011 : out <= 16'sb11111111_10101110; // -0.32241
        11'b10001101100 : out <= 16'sb11111111_10101101; // -0.32531
        11'b10001101101 : out <= 16'sb11111111_10101100; // -0.32821
        11'b10001101110 : out <= 16'sb11111111_10101100; // -0.33111
        11'b10001101111 : out <= 16'sb11111111_10101011; // -0.33400
        11'b10001110000 : out <= 16'sb11111111_10101010; // -0.33689
        11'b10001110001 : out <= 16'sb11111111_10101010; // -0.33978
        11'b10001110010 : out <= 16'sb11111111_10101001; // -0.34266
        11'b10001110011 : out <= 16'sb11111111_10101000; // -0.34554
        11'b10001110100 : out <= 16'sb11111111_10100111; // -0.34842
        11'b10001110101 : out <= 16'sb11111111_10100111; // -0.35129
        11'b10001110110 : out <= 16'sb11111111_10100110; // -0.35416
        11'b10001110111 : out <= 16'sb11111111_10100101; // -0.35703
        11'b10001111000 : out <= 16'sb11111111_10100100; // -0.35990
        11'b10001111001 : out <= 16'sb11111111_10100100; // -0.36276
        11'b10001111010 : out <= 16'sb11111111_10100011; // -0.36561
        11'b10001111011 : out <= 16'sb11111111_10100010; // -0.36847
        11'b10001111100 : out <= 16'sb11111111_10100001; // -0.37132
        11'b10001111101 : out <= 16'sb11111111_10100001; // -0.37416
        11'b10001111110 : out <= 16'sb11111111_10100000; // -0.37701
        11'b10001111111 : out <= 16'sb11111111_10011111; // -0.37985
        11'b10010000000 : out <= 16'sb11111111_10011111; // -0.38268
        11'b10010000001 : out <= 16'sb11111111_10011110; // -0.38552
        11'b10010000010 : out <= 16'sb11111111_10011101; // -0.38835
        11'b10010000011 : out <= 16'sb11111111_10011100; // -0.39117
        11'b10010000100 : out <= 16'sb11111111_10011100; // -0.39399
        11'b10010000101 : out <= 16'sb11111111_10011011; // -0.39681
        11'b10010000110 : out <= 16'sb11111111_10011010; // -0.39962
        11'b10010000111 : out <= 16'sb11111111_10011001; // -0.40243
        11'b10010001000 : out <= 16'sb11111111_10011001; // -0.40524
        11'b10010001001 : out <= 16'sb11111111_10011000; // -0.40804
        11'b10010001010 : out <= 16'sb11111111_10010111; // -0.41084
        11'b10010001011 : out <= 16'sb11111111_10010111; // -0.41364
        11'b10010001100 : out <= 16'sb11111111_10010110; // -0.41643
        11'b10010001101 : out <= 16'sb11111111_10010101; // -0.41922
        11'b10010001110 : out <= 16'sb11111111_10010100; // -0.42200
        11'b10010001111 : out <= 16'sb11111111_10010100; // -0.42478
        11'b10010010000 : out <= 16'sb11111111_10010011; // -0.42756
        11'b10010010001 : out <= 16'sb11111111_10010010; // -0.43033
        11'b10010010010 : out <= 16'sb11111111_10010010; // -0.43309
        11'b10010010011 : out <= 16'sb11111111_10010001; // -0.43586
        11'b10010010100 : out <= 16'sb11111111_10010000; // -0.43862
        11'b10010010101 : out <= 16'sb11111111_10010000; // -0.44137
        11'b10010010110 : out <= 16'sb11111111_10001111; // -0.44412
        11'b10010010111 : out <= 16'sb11111111_10001110; // -0.44687
        11'b10010011000 : out <= 16'sb11111111_10001101; // -0.44961
        11'b10010011001 : out <= 16'sb11111111_10001101; // -0.45235
        11'b10010011010 : out <= 16'sb11111111_10001100; // -0.45508
        11'b10010011011 : out <= 16'sb11111111_10001011; // -0.45781
        11'b10010011100 : out <= 16'sb11111111_10001011; // -0.46054
        11'b10010011101 : out <= 16'sb11111111_10001010; // -0.46326
        11'b10010011110 : out <= 16'sb11111111_10001001; // -0.46598
        11'b10010011111 : out <= 16'sb11111111_10001001; // -0.46869
        11'b10010100000 : out <= 16'sb11111111_10001000; // -0.47140
        11'b10010100001 : out <= 16'sb11111111_10000111; // -0.47410
        11'b10010100010 : out <= 16'sb11111111_10000110; // -0.47680
        11'b10010100011 : out <= 16'sb11111111_10000110; // -0.47949
        11'b10010100100 : out <= 16'sb11111111_10000101; // -0.48218
        11'b10010100101 : out <= 16'sb11111111_10000100; // -0.48487
        11'b10010100110 : out <= 16'sb11111111_10000100; // -0.48755
        11'b10010100111 : out <= 16'sb11111111_10000011; // -0.49023
        11'b10010101000 : out <= 16'sb11111111_10000010; // -0.49290
        11'b10010101001 : out <= 16'sb11111111_10000010; // -0.49557
        11'b10010101010 : out <= 16'sb11111111_10000001; // -0.49823
        11'b10010101011 : out <= 16'sb11111111_10000000; // -0.50089
        11'b10010101100 : out <= 16'sb11111111_10000000; // -0.50354
        11'b10010101101 : out <= 16'sb11111111_01111111; // -0.50619
        11'b10010101110 : out <= 16'sb11111111_01111110; // -0.50883
        11'b10010101111 : out <= 16'sb11111111_01111110; // -0.51147
        11'b10010110000 : out <= 16'sb11111111_01111101; // -0.51410
        11'b10010110001 : out <= 16'sb11111111_01111100; // -0.51673
        11'b10010110010 : out <= 16'sb11111111_01111100; // -0.51936
        11'b10010110011 : out <= 16'sb11111111_01111011; // -0.52198
        11'b10010110100 : out <= 16'sb11111111_01111010; // -0.52459
        11'b10010110101 : out <= 16'sb11111111_01111010; // -0.52720
        11'b10010110110 : out <= 16'sb11111111_01111001; // -0.52980
        11'b10010110111 : out <= 16'sb11111111_01111000; // -0.53240
        11'b10010111000 : out <= 16'sb11111111_01111000; // -0.53500
        11'b10010111001 : out <= 16'sb11111111_01110111; // -0.53759
        11'b10010111010 : out <= 16'sb11111111_01110110; // -0.54017
        11'b10010111011 : out <= 16'sb11111111_01110110; // -0.54275
        11'b10010111100 : out <= 16'sb11111111_01110101; // -0.54532
        11'b10010111101 : out <= 16'sb11111111_01110100; // -0.54789
        11'b10010111110 : out <= 16'sb11111111_01110100; // -0.55046
        11'b10010111111 : out <= 16'sb11111111_01110011; // -0.55302
        11'b10011000000 : out <= 16'sb11111111_01110010; // -0.55557
        11'b10011000001 : out <= 16'sb11111111_01110010; // -0.55812
        11'b10011000010 : out <= 16'sb11111111_01110001; // -0.56066
        11'b10011000011 : out <= 16'sb11111111_01110000; // -0.56320
        11'b10011000100 : out <= 16'sb11111111_01110000; // -0.56573
        11'b10011000101 : out <= 16'sb11111111_01101111; // -0.56826
        11'b10011000110 : out <= 16'sb11111111_01101110; // -0.57078
        11'b10011000111 : out <= 16'sb11111111_01101110; // -0.57330
        11'b10011001000 : out <= 16'sb11111111_01101101; // -0.57581
        11'b10011001001 : out <= 16'sb11111111_01101100; // -0.57831
        11'b10011001010 : out <= 16'sb11111111_01101100; // -0.58081
        11'b10011001011 : out <= 16'sb11111111_01101011; // -0.58331
        11'b10011001100 : out <= 16'sb11111111_01101011; // -0.58580
        11'b10011001101 : out <= 16'sb11111111_01101010; // -0.58828
        11'b10011001110 : out <= 16'sb11111111_01101001; // -0.59076
        11'b10011001111 : out <= 16'sb11111111_01101001; // -0.59323
        11'b10011010000 : out <= 16'sb11111111_01101000; // -0.59570
        11'b10011010001 : out <= 16'sb11111111_01100111; // -0.59816
        11'b10011010010 : out <= 16'sb11111111_01100111; // -0.60062
        11'b10011010011 : out <= 16'sb11111111_01100110; // -0.60307
        11'b10011010100 : out <= 16'sb11111111_01100101; // -0.60551
        11'b10011010101 : out <= 16'sb11111111_01100101; // -0.60795
        11'b10011010110 : out <= 16'sb11111111_01100100; // -0.61038
        11'b10011010111 : out <= 16'sb11111111_01100100; // -0.61281
        11'b10011011000 : out <= 16'sb11111111_01100011; // -0.61523
        11'b10011011001 : out <= 16'sb11111111_01100010; // -0.61765
        11'b10011011010 : out <= 16'sb11111111_01100010; // -0.62006
        11'b10011011011 : out <= 16'sb11111111_01100001; // -0.62246
        11'b10011011100 : out <= 16'sb11111111_01100001; // -0.62486
        11'b10011011101 : out <= 16'sb11111111_01100000; // -0.62725
        11'b10011011110 : out <= 16'sb11111111_01011111; // -0.62964
        11'b10011011111 : out <= 16'sb11111111_01011111; // -0.63202
        11'b10011100000 : out <= 16'sb11111111_01011110; // -0.63439
        11'b10011100001 : out <= 16'sb11111111_01011101; // -0.63676
        11'b10011100010 : out <= 16'sb11111111_01011101; // -0.63912
        11'b10011100011 : out <= 16'sb11111111_01011100; // -0.64148
        11'b10011100100 : out <= 16'sb11111111_01011100; // -0.64383
        11'b10011100101 : out <= 16'sb11111111_01011011; // -0.64618
        11'b10011100110 : out <= 16'sb11111111_01011010; // -0.64851
        11'b10011100111 : out <= 16'sb11111111_01011010; // -0.65085
        11'b10011101000 : out <= 16'sb11111111_01011001; // -0.65317
        11'b10011101001 : out <= 16'sb11111111_01011001; // -0.65549
        11'b10011101010 : out <= 16'sb11111111_01011000; // -0.65781
        11'b10011101011 : out <= 16'sb11111111_01011000; // -0.66011
        11'b10011101100 : out <= 16'sb11111111_01010111; // -0.66242
        11'b10011101101 : out <= 16'sb11111111_01010110; // -0.66471
        11'b10011101110 : out <= 16'sb11111111_01010110; // -0.66700
        11'b10011101111 : out <= 16'sb11111111_01010101; // -0.66928
        11'b10011110000 : out <= 16'sb11111111_01010101; // -0.67156
        11'b10011110001 : out <= 16'sb11111111_01010100; // -0.67383
        11'b10011110010 : out <= 16'sb11111111_01010011; // -0.67609
        11'b10011110011 : out <= 16'sb11111111_01010011; // -0.67835
        11'b10011110100 : out <= 16'sb11111111_01010010; // -0.68060
        11'b10011110101 : out <= 16'sb11111111_01010010; // -0.68285
        11'b10011110110 : out <= 16'sb11111111_01010001; // -0.68508
        11'b10011110111 : out <= 16'sb11111111_01010001; // -0.68732
        11'b10011111000 : out <= 16'sb11111111_01010000; // -0.68954
        11'b10011111001 : out <= 16'sb11111111_01001111; // -0.69176
        11'b10011111010 : out <= 16'sb11111111_01001111; // -0.69397
        11'b10011111011 : out <= 16'sb11111111_01001110; // -0.69618
        11'b10011111100 : out <= 16'sb11111111_01001110; // -0.69838
        11'b10011111101 : out <= 16'sb11111111_01001101; // -0.70057
        11'b10011111110 : out <= 16'sb11111111_01001101; // -0.70275
        11'b10011111111 : out <= 16'sb11111111_01001100; // -0.70493
        11'b10100000000 : out <= 16'sb11111111_01001011; // -0.70711
        11'b10100000001 : out <= 16'sb11111111_01001011; // -0.70927
        11'b10100000010 : out <= 16'sb11111111_01001010; // -0.71143
        11'b10100000011 : out <= 16'sb11111111_01001010; // -0.71358
        11'b10100000100 : out <= 16'sb11111111_01001001; // -0.71573
        11'b10100000101 : out <= 16'sb11111111_01001001; // -0.71787
        11'b10100000110 : out <= 16'sb11111111_01001000; // -0.72000
        11'b10100000111 : out <= 16'sb11111111_01001000; // -0.72213
        11'b10100001000 : out <= 16'sb11111111_01000111; // -0.72425
        11'b10100001001 : out <= 16'sb11111111_01000111; // -0.72636
        11'b10100001010 : out <= 16'sb11111111_01000110; // -0.72846
        11'b10100001011 : out <= 16'sb11111111_01000101; // -0.73056
        11'b10100001100 : out <= 16'sb11111111_01000101; // -0.73265
        11'b10100001101 : out <= 16'sb11111111_01000100; // -0.73474
        11'b10100001110 : out <= 16'sb11111111_01000100; // -0.73682
        11'b10100001111 : out <= 16'sb11111111_01000011; // -0.73889
        11'b10100010000 : out <= 16'sb11111111_01000011; // -0.74095
        11'b10100010001 : out <= 16'sb11111111_01000010; // -0.74301
        11'b10100010010 : out <= 16'sb11111111_01000010; // -0.74506
        11'b10100010011 : out <= 16'sb11111111_01000001; // -0.74710
        11'b10100010100 : out <= 16'sb11111111_01000001; // -0.74914
        11'b10100010101 : out <= 16'sb11111111_01000000; // -0.75117
        11'b10100010110 : out <= 16'sb11111111_01000000; // -0.75319
        11'b10100010111 : out <= 16'sb11111111_00111111; // -0.75520
        11'b10100011000 : out <= 16'sb11111111_00111111; // -0.75721
        11'b10100011001 : out <= 16'sb11111111_00111110; // -0.75921
        11'b10100011010 : out <= 16'sb11111111_00111110; // -0.76120
        11'b10100011011 : out <= 16'sb11111111_00111101; // -0.76319
        11'b10100011100 : out <= 16'sb11111111_00111101; // -0.76517
        11'b10100011101 : out <= 16'sb11111111_00111100; // -0.76714
        11'b10100011110 : out <= 16'sb11111111_00111100; // -0.76910
        11'b10100011111 : out <= 16'sb11111111_00111011; // -0.77106
        11'b10100100000 : out <= 16'sb11111111_00111011; // -0.77301
        11'b10100100001 : out <= 16'sb11111111_00111010; // -0.77495
        11'b10100100010 : out <= 16'sb11111111_00111010; // -0.77689
        11'b10100100011 : out <= 16'sb11111111_00111001; // -0.77882
        11'b10100100100 : out <= 16'sb11111111_00111001; // -0.78074
        11'b10100100101 : out <= 16'sb11111111_00111000; // -0.78265
        11'b10100100110 : out <= 16'sb11111111_00111000; // -0.78456
        11'b10100100111 : out <= 16'sb11111111_00110111; // -0.78646
        11'b10100101000 : out <= 16'sb11111111_00110111; // -0.78835
        11'b10100101001 : out <= 16'sb11111111_00110110; // -0.79023
        11'b10100101010 : out <= 16'sb11111111_00110110; // -0.79211
        11'b10100101011 : out <= 16'sb11111111_00110101; // -0.79398
        11'b10100101100 : out <= 16'sb11111111_00110101; // -0.79584
        11'b10100101101 : out <= 16'sb11111111_00110100; // -0.79769
        11'b10100101110 : out <= 16'sb11111111_00110100; // -0.79954
        11'b10100101111 : out <= 16'sb11111111_00110011; // -0.80138
        11'b10100110000 : out <= 16'sb11111111_00110011; // -0.80321
        11'b10100110001 : out <= 16'sb11111111_00110010; // -0.80503
        11'b10100110010 : out <= 16'sb11111111_00110010; // -0.80685
        11'b10100110011 : out <= 16'sb11111111_00110001; // -0.80866
        11'b10100110100 : out <= 16'sb11111111_00110001; // -0.81046
        11'b10100110101 : out <= 16'sb11111111_00110001; // -0.81225
        11'b10100110110 : out <= 16'sb11111111_00110000; // -0.81404
        11'b10100110111 : out <= 16'sb11111111_00110000; // -0.81581
        11'b10100111000 : out <= 16'sb11111111_00101111; // -0.81758
        11'b10100111001 : out <= 16'sb11111111_00101111; // -0.81935
        11'b10100111010 : out <= 16'sb11111111_00101110; // -0.82110
        11'b10100111011 : out <= 16'sb11111111_00101110; // -0.82285
        11'b10100111100 : out <= 16'sb11111111_00101101; // -0.82459
        11'b10100111101 : out <= 16'sb11111111_00101101; // -0.82632
        11'b10100111110 : out <= 16'sb11111111_00101101; // -0.82805
        11'b10100111111 : out <= 16'sb11111111_00101100; // -0.82976
        11'b10101000000 : out <= 16'sb11111111_00101100; // -0.83147
        11'b10101000001 : out <= 16'sb11111111_00101011; // -0.83317
        11'b10101000010 : out <= 16'sb11111111_00101011; // -0.83486
        11'b10101000011 : out <= 16'sb11111111_00101010; // -0.83655
        11'b10101000100 : out <= 16'sb11111111_00101010; // -0.83822
        11'b10101000101 : out <= 16'sb11111111_00101001; // -0.83989
        11'b10101000110 : out <= 16'sb11111111_00101001; // -0.84155
        11'b10101000111 : out <= 16'sb11111111_00101001; // -0.84321
        11'b10101001000 : out <= 16'sb11111111_00101000; // -0.84485
        11'b10101001001 : out <= 16'sb11111111_00101000; // -0.84649
        11'b10101001010 : out <= 16'sb11111111_00100111; // -0.84812
        11'b10101001011 : out <= 16'sb11111111_00100111; // -0.84974
        11'b10101001100 : out <= 16'sb11111111_00100111; // -0.85136
        11'b10101001101 : out <= 16'sb11111111_00100110; // -0.85296
        11'b10101001110 : out <= 16'sb11111111_00100110; // -0.85456
        11'b10101001111 : out <= 16'sb11111111_00100101; // -0.85615
        11'b10101010000 : out <= 16'sb11111111_00100101; // -0.85773
        11'b10101010001 : out <= 16'sb11111111_00100101; // -0.85930
        11'b10101010010 : out <= 16'sb11111111_00100100; // -0.86087
        11'b10101010011 : out <= 16'sb11111111_00100100; // -0.86242
        11'b10101010100 : out <= 16'sb11111111_00100011; // -0.86397
        11'b10101010101 : out <= 16'sb11111111_00100011; // -0.86551
        11'b10101010110 : out <= 16'sb11111111_00100011; // -0.86705
        11'b10101010111 : out <= 16'sb11111111_00100010; // -0.86857
        11'b10101011000 : out <= 16'sb11111111_00100010; // -0.87009
        11'b10101011001 : out <= 16'sb11111111_00100001; // -0.87160
        11'b10101011010 : out <= 16'sb11111111_00100001; // -0.87309
        11'b10101011011 : out <= 16'sb11111111_00100001; // -0.87459
        11'b10101011100 : out <= 16'sb11111111_00100000; // -0.87607
        11'b10101011101 : out <= 16'sb11111111_00100000; // -0.87755
        11'b10101011110 : out <= 16'sb11111111_00011111; // -0.87901
        11'b10101011111 : out <= 16'sb11111111_00011111; // -0.88047
        11'b10101100000 : out <= 16'sb11111111_00011111; // -0.88192
        11'b10101100001 : out <= 16'sb11111111_00011110; // -0.88336
        11'b10101100010 : out <= 16'sb11111111_00011110; // -0.88480
        11'b10101100011 : out <= 16'sb11111111_00011110; // -0.88622
        11'b10101100100 : out <= 16'sb11111111_00011101; // -0.88764
        11'b10101100101 : out <= 16'sb11111111_00011101; // -0.88905
        11'b10101100110 : out <= 16'sb11111111_00011101; // -0.89045
        11'b10101100111 : out <= 16'sb11111111_00011100; // -0.89184
        11'b10101101000 : out <= 16'sb11111111_00011100; // -0.89322
        11'b10101101001 : out <= 16'sb11111111_00011011; // -0.89460
        11'b10101101010 : out <= 16'sb11111111_00011011; // -0.89597
        11'b10101101011 : out <= 16'sb11111111_00011011; // -0.89732
        11'b10101101100 : out <= 16'sb11111111_00011010; // -0.89867
        11'b10101101101 : out <= 16'sb11111111_00011010; // -0.90002
        11'b10101101110 : out <= 16'sb11111111_00011010; // -0.90135
        11'b10101101111 : out <= 16'sb11111111_00011001; // -0.90267
        11'b10101110000 : out <= 16'sb11111111_00011001; // -0.90399
        11'b10101110001 : out <= 16'sb11111111_00011001; // -0.90530
        11'b10101110010 : out <= 16'sb11111111_00011000; // -0.90660
        11'b10101110011 : out <= 16'sb11111111_00011000; // -0.90789
        11'b10101110100 : out <= 16'sb11111111_00011000; // -0.90917
        11'b10101110101 : out <= 16'sb11111111_00010111; // -0.91044
        11'b10101110110 : out <= 16'sb11111111_00010111; // -0.91171
        11'b10101110111 : out <= 16'sb11111111_00010111; // -0.91296
        11'b10101111000 : out <= 16'sb11111111_00010110; // -0.91421
        11'b10101111001 : out <= 16'sb11111111_00010110; // -0.91545
        11'b10101111010 : out <= 16'sb11111111_00010110; // -0.91668
        11'b10101111011 : out <= 16'sb11111111_00010110; // -0.91790
        11'b10101111100 : out <= 16'sb11111111_00010101; // -0.91911
        11'b10101111101 : out <= 16'sb11111111_00010101; // -0.92032
        11'b10101111110 : out <= 16'sb11111111_00010101; // -0.92151
        11'b10101111111 : out <= 16'sb11111111_00010100; // -0.92270
        11'b10110000000 : out <= 16'sb11111111_00010100; // -0.92388
        11'b10110000001 : out <= 16'sb11111111_00010100; // -0.92505
        11'b10110000010 : out <= 16'sb11111111_00010011; // -0.92621
        11'b10110000011 : out <= 16'sb11111111_00010011; // -0.92736
        11'b10110000100 : out <= 16'sb11111111_00010011; // -0.92851
        11'b10110000101 : out <= 16'sb11111111_00010011; // -0.92964
        11'b10110000110 : out <= 16'sb11111111_00010010; // -0.93077
        11'b10110000111 : out <= 16'sb11111111_00010010; // -0.93188
        11'b10110001000 : out <= 16'sb11111111_00010010; // -0.93299
        11'b10110001001 : out <= 16'sb11111111_00010001; // -0.93409
        11'b10110001010 : out <= 16'sb11111111_00010001; // -0.93518
        11'b10110001011 : out <= 16'sb11111111_00010001; // -0.93627
        11'b10110001100 : out <= 16'sb11111111_00010001; // -0.93734
        11'b10110001101 : out <= 16'sb11111111_00010000; // -0.93840
        11'b10110001110 : out <= 16'sb11111111_00010000; // -0.93946
        11'b10110001111 : out <= 16'sb11111111_00010000; // -0.94051
        11'b10110010000 : out <= 16'sb11111111_00001111; // -0.94154
        11'b10110010001 : out <= 16'sb11111111_00001111; // -0.94257
        11'b10110010010 : out <= 16'sb11111111_00001111; // -0.94359
        11'b10110010011 : out <= 16'sb11111111_00001111; // -0.94460
        11'b10110010100 : out <= 16'sb11111111_00001110; // -0.94561
        11'b10110010101 : out <= 16'sb11111111_00001110; // -0.94660
        11'b10110010110 : out <= 16'sb11111111_00001110; // -0.94759
        11'b10110010111 : out <= 16'sb11111111_00001110; // -0.94856
        11'b10110011000 : out <= 16'sb11111111_00001101; // -0.94953
        11'b10110011001 : out <= 16'sb11111111_00001101; // -0.95049
        11'b10110011010 : out <= 16'sb11111111_00001101; // -0.95144
        11'b10110011011 : out <= 16'sb11111111_00001101; // -0.95238
        11'b10110011100 : out <= 16'sb11111111_00001100; // -0.95331
        11'b10110011101 : out <= 16'sb11111111_00001100; // -0.95423
        11'b10110011110 : out <= 16'sb11111111_00001100; // -0.95514
        11'b10110011111 : out <= 16'sb11111111_00001100; // -0.95605
        11'b10110100000 : out <= 16'sb11111111_00001100; // -0.95694
        11'b10110100001 : out <= 16'sb11111111_00001011; // -0.95783
        11'b10110100010 : out <= 16'sb11111111_00001011; // -0.95870
        11'b10110100011 : out <= 16'sb11111111_00001011; // -0.95957
        11'b10110100100 : out <= 16'sb11111111_00001011; // -0.96043
        11'b10110100101 : out <= 16'sb11111111_00001010; // -0.96128
        11'b10110100110 : out <= 16'sb11111111_00001010; // -0.96212
        11'b10110100111 : out <= 16'sb11111111_00001010; // -0.96295
        11'b10110101000 : out <= 16'sb11111111_00001010; // -0.96378
        11'b10110101001 : out <= 16'sb11111111_00001010; // -0.96459
        11'b10110101010 : out <= 16'sb11111111_00001001; // -0.96539
        11'b10110101011 : out <= 16'sb11111111_00001001; // -0.96619
        11'b10110101100 : out <= 16'sb11111111_00001001; // -0.96698
        11'b10110101101 : out <= 16'sb11111111_00001001; // -0.96775
        11'b10110101110 : out <= 16'sb11111111_00001001; // -0.96852
        11'b10110101111 : out <= 16'sb11111111_00001000; // -0.96928
        11'b10110110000 : out <= 16'sb11111111_00001000; // -0.97003
        11'b10110110001 : out <= 16'sb11111111_00001000; // -0.97077
        11'b10110110010 : out <= 16'sb11111111_00001000; // -0.97150
        11'b10110110011 : out <= 16'sb11111111_00001000; // -0.97223
        11'b10110110100 : out <= 16'sb11111111_00000111; // -0.97294
        11'b10110110101 : out <= 16'sb11111111_00000111; // -0.97364
        11'b10110110110 : out <= 16'sb11111111_00000111; // -0.97434
        11'b10110110111 : out <= 16'sb11111111_00000111; // -0.97503
        11'b10110111000 : out <= 16'sb11111111_00000111; // -0.97570
        11'b10110111001 : out <= 16'sb11111111_00000111; // -0.97637
        11'b10110111010 : out <= 16'sb11111111_00000110; // -0.97703
        11'b10110111011 : out <= 16'sb11111111_00000110; // -0.97768
        11'b10110111100 : out <= 16'sb11111111_00000110; // -0.97832
        11'b10110111101 : out <= 16'sb11111111_00000110; // -0.97895
        11'b10110111110 : out <= 16'sb11111111_00000110; // -0.97957
        11'b10110111111 : out <= 16'sb11111111_00000110; // -0.98018
        11'b10111000000 : out <= 16'sb11111111_00000101; // -0.98079
        11'b10111000001 : out <= 16'sb11111111_00000101; // -0.98138
        11'b10111000010 : out <= 16'sb11111111_00000101; // -0.98196
        11'b10111000011 : out <= 16'sb11111111_00000101; // -0.98254
        11'b10111000100 : out <= 16'sb11111111_00000101; // -0.98311
        11'b10111000101 : out <= 16'sb11111111_00000101; // -0.98366
        11'b10111000110 : out <= 16'sb11111111_00000101; // -0.98421
        11'b10111000111 : out <= 16'sb11111111_00000100; // -0.98475
        11'b10111001000 : out <= 16'sb11111111_00000100; // -0.98528
        11'b10111001001 : out <= 16'sb11111111_00000100; // -0.98580
        11'b10111001010 : out <= 16'sb11111111_00000100; // -0.98631
        11'b10111001011 : out <= 16'sb11111111_00000100; // -0.98681
        11'b10111001100 : out <= 16'sb11111111_00000100; // -0.98730
        11'b10111001101 : out <= 16'sb11111111_00000100; // -0.98778
        11'b10111001110 : out <= 16'sb11111111_00000100; // -0.98826
        11'b10111001111 : out <= 16'sb11111111_00000011; // -0.98872
        11'b10111010000 : out <= 16'sb11111111_00000011; // -0.98918
        11'b10111010001 : out <= 16'sb11111111_00000011; // -0.98962
        11'b10111010010 : out <= 16'sb11111111_00000011; // -0.99006
        11'b10111010011 : out <= 16'sb11111111_00000011; // -0.99049
        11'b10111010100 : out <= 16'sb11111111_00000011; // -0.99090
        11'b10111010101 : out <= 16'sb11111111_00000011; // -0.99131
        11'b10111010110 : out <= 16'sb11111111_00000011; // -0.99171
        11'b10111010111 : out <= 16'sb11111111_00000011; // -0.99210
        11'b10111011000 : out <= 16'sb11111111_00000010; // -0.99248
        11'b10111011001 : out <= 16'sb11111111_00000010; // -0.99285
        11'b10111011010 : out <= 16'sb11111111_00000010; // -0.99321
        11'b10111011011 : out <= 16'sb11111111_00000010; // -0.99356
        11'b10111011100 : out <= 16'sb11111111_00000010; // -0.99391
        11'b10111011101 : out <= 16'sb11111111_00000010; // -0.99424
        11'b10111011110 : out <= 16'sb11111111_00000010; // -0.99456
        11'b10111011111 : out <= 16'sb11111111_00000010; // -0.99488
        11'b10111100000 : out <= 16'sb11111111_00000010; // -0.99518
        11'b10111100001 : out <= 16'sb11111111_00000010; // -0.99548
        11'b10111100010 : out <= 16'sb11111111_00000010; // -0.99577
        11'b10111100011 : out <= 16'sb11111111_00000010; // -0.99604
        11'b10111100100 : out <= 16'sb11111111_00000001; // -0.99631
        11'b10111100101 : out <= 16'sb11111111_00000001; // -0.99657
        11'b10111100110 : out <= 16'sb11111111_00000001; // -0.99682
        11'b10111100111 : out <= 16'sb11111111_00000001; // -0.99706
        11'b10111101000 : out <= 16'sb11111111_00000001; // -0.99729
        11'b10111101001 : out <= 16'sb11111111_00000001; // -0.99751
        11'b10111101010 : out <= 16'sb11111111_00000001; // -0.99772
        11'b10111101011 : out <= 16'sb11111111_00000001; // -0.99793
        11'b10111101100 : out <= 16'sb11111111_00000001; // -0.99812
        11'b10111101101 : out <= 16'sb11111111_00000001; // -0.99830
        11'b10111101110 : out <= 16'sb11111111_00000001; // -0.99848
        11'b10111101111 : out <= 16'sb11111111_00000001; // -0.99864
        11'b10111110000 : out <= 16'sb11111111_00000001; // -0.99880
        11'b10111110001 : out <= 16'sb11111111_00000001; // -0.99894
        11'b10111110010 : out <= 16'sb11111111_00000001; // -0.99908
        11'b10111110011 : out <= 16'sb11111111_00000001; // -0.99920
        11'b10111110100 : out <= 16'sb11111111_00000001; // -0.99932
        11'b10111110101 : out <= 16'sb11111111_00000001; // -0.99943
        11'b10111110110 : out <= 16'sb11111111_00000001; // -0.99953
        11'b10111110111 : out <= 16'sb11111111_00000001; // -0.99962
        11'b10111111000 : out <= 16'sb11111111_00000001; // -0.99970
        11'b10111111001 : out <= 16'sb11111111_00000001; // -0.99977
        11'b10111111010 : out <= 16'sb11111111_00000001; // -0.99983
        11'b10111111011 : out <= 16'sb11111111_00000001; // -0.99988
        11'b10111111100 : out <= 16'sb11111111_00000001; // -0.99992
        11'b10111111101 : out <= 16'sb11111111_00000001; // -0.99996
        11'b10111111110 : out <= 16'sb11111111_00000001; // -0.99998
        11'b10111111111 : out <= 16'sb11111111_00000001; // -1.00000
        11'b11000000000 : out <= 16'sb11111111_00000000; // -1.00000
        11'b11000000001 : out <= 16'sb11111111_00000001; // -1.00000
        11'b11000000010 : out <= 16'sb11111111_00000001; // -0.99998
        11'b11000000011 : out <= 16'sb11111111_00000001; // -0.99996
        11'b11000000100 : out <= 16'sb11111111_00000001; // -0.99992
        11'b11000000101 : out <= 16'sb11111111_00000001; // -0.99988
        11'b11000000110 : out <= 16'sb11111111_00000001; // -0.99983
        11'b11000000111 : out <= 16'sb11111111_00000001; // -0.99977
        11'b11000001000 : out <= 16'sb11111111_00000001; // -0.99970
        11'b11000001001 : out <= 16'sb11111111_00000001; // -0.99962
        11'b11000001010 : out <= 16'sb11111111_00000001; // -0.99953
        11'b11000001011 : out <= 16'sb11111111_00000001; // -0.99943
        11'b11000001100 : out <= 16'sb11111111_00000001; // -0.99932
        11'b11000001101 : out <= 16'sb11111111_00000001; // -0.99920
        11'b11000001110 : out <= 16'sb11111111_00000001; // -0.99908
        11'b11000001111 : out <= 16'sb11111111_00000001; // -0.99894
        11'b11000010000 : out <= 16'sb11111111_00000001; // -0.99880
        11'b11000010001 : out <= 16'sb11111111_00000001; // -0.99864
        11'b11000010010 : out <= 16'sb11111111_00000001; // -0.99848
        11'b11000010011 : out <= 16'sb11111111_00000001; // -0.99830
        11'b11000010100 : out <= 16'sb11111111_00000001; // -0.99812
        11'b11000010101 : out <= 16'sb11111111_00000001; // -0.99793
        11'b11000010110 : out <= 16'sb11111111_00000001; // -0.99772
        11'b11000010111 : out <= 16'sb11111111_00000001; // -0.99751
        11'b11000011000 : out <= 16'sb11111111_00000001; // -0.99729
        11'b11000011001 : out <= 16'sb11111111_00000001; // -0.99706
        11'b11000011010 : out <= 16'sb11111111_00000001; // -0.99682
        11'b11000011011 : out <= 16'sb11111111_00000001; // -0.99657
        11'b11000011100 : out <= 16'sb11111111_00000001; // -0.99631
        11'b11000011101 : out <= 16'sb11111111_00000010; // -0.99604
        11'b11000011110 : out <= 16'sb11111111_00000010; // -0.99577
        11'b11000011111 : out <= 16'sb11111111_00000010; // -0.99548
        11'b11000100000 : out <= 16'sb11111111_00000010; // -0.99518
        11'b11000100001 : out <= 16'sb11111111_00000010; // -0.99488
        11'b11000100010 : out <= 16'sb11111111_00000010; // -0.99456
        11'b11000100011 : out <= 16'sb11111111_00000010; // -0.99424
        11'b11000100100 : out <= 16'sb11111111_00000010; // -0.99391
        11'b11000100101 : out <= 16'sb11111111_00000010; // -0.99356
        11'b11000100110 : out <= 16'sb11111111_00000010; // -0.99321
        11'b11000100111 : out <= 16'sb11111111_00000010; // -0.99285
        11'b11000101000 : out <= 16'sb11111111_00000010; // -0.99248
        11'b11000101001 : out <= 16'sb11111111_00000011; // -0.99210
        11'b11000101010 : out <= 16'sb11111111_00000011; // -0.99171
        11'b11000101011 : out <= 16'sb11111111_00000011; // -0.99131
        11'b11000101100 : out <= 16'sb11111111_00000011; // -0.99090
        11'b11000101101 : out <= 16'sb11111111_00000011; // -0.99049
        11'b11000101110 : out <= 16'sb11111111_00000011; // -0.99006
        11'b11000101111 : out <= 16'sb11111111_00000011; // -0.98962
        11'b11000110000 : out <= 16'sb11111111_00000011; // -0.98918
        11'b11000110001 : out <= 16'sb11111111_00000011; // -0.98872
        11'b11000110010 : out <= 16'sb11111111_00000100; // -0.98826
        11'b11000110011 : out <= 16'sb11111111_00000100; // -0.98778
        11'b11000110100 : out <= 16'sb11111111_00000100; // -0.98730
        11'b11000110101 : out <= 16'sb11111111_00000100; // -0.98681
        11'b11000110110 : out <= 16'sb11111111_00000100; // -0.98631
        11'b11000110111 : out <= 16'sb11111111_00000100; // -0.98580
        11'b11000111000 : out <= 16'sb11111111_00000100; // -0.98528
        11'b11000111001 : out <= 16'sb11111111_00000100; // -0.98475
        11'b11000111010 : out <= 16'sb11111111_00000101; // -0.98421
        11'b11000111011 : out <= 16'sb11111111_00000101; // -0.98366
        11'b11000111100 : out <= 16'sb11111111_00000101; // -0.98311
        11'b11000111101 : out <= 16'sb11111111_00000101; // -0.98254
        11'b11000111110 : out <= 16'sb11111111_00000101; // -0.98196
        11'b11000111111 : out <= 16'sb11111111_00000101; // -0.98138
        11'b11001000000 : out <= 16'sb11111111_00000101; // -0.98079
        11'b11001000001 : out <= 16'sb11111111_00000110; // -0.98018
        11'b11001000010 : out <= 16'sb11111111_00000110; // -0.97957
        11'b11001000011 : out <= 16'sb11111111_00000110; // -0.97895
        11'b11001000100 : out <= 16'sb11111111_00000110; // -0.97832
        11'b11001000101 : out <= 16'sb11111111_00000110; // -0.97768
        11'b11001000110 : out <= 16'sb11111111_00000110; // -0.97703
        11'b11001000111 : out <= 16'sb11111111_00000111; // -0.97637
        11'b11001001000 : out <= 16'sb11111111_00000111; // -0.97570
        11'b11001001001 : out <= 16'sb11111111_00000111; // -0.97503
        11'b11001001010 : out <= 16'sb11111111_00000111; // -0.97434
        11'b11001001011 : out <= 16'sb11111111_00000111; // -0.97364
        11'b11001001100 : out <= 16'sb11111111_00000111; // -0.97294
        11'b11001001101 : out <= 16'sb11111111_00001000; // -0.97223
        11'b11001001110 : out <= 16'sb11111111_00001000; // -0.97150
        11'b11001001111 : out <= 16'sb11111111_00001000; // -0.97077
        11'b11001010000 : out <= 16'sb11111111_00001000; // -0.97003
        11'b11001010001 : out <= 16'sb11111111_00001000; // -0.96928
        11'b11001010010 : out <= 16'sb11111111_00001001; // -0.96852
        11'b11001010011 : out <= 16'sb11111111_00001001; // -0.96775
        11'b11001010100 : out <= 16'sb11111111_00001001; // -0.96698
        11'b11001010101 : out <= 16'sb11111111_00001001; // -0.96619
        11'b11001010110 : out <= 16'sb11111111_00001001; // -0.96539
        11'b11001010111 : out <= 16'sb11111111_00001010; // -0.96459
        11'b11001011000 : out <= 16'sb11111111_00001010; // -0.96378
        11'b11001011001 : out <= 16'sb11111111_00001010; // -0.96295
        11'b11001011010 : out <= 16'sb11111111_00001010; // -0.96212
        11'b11001011011 : out <= 16'sb11111111_00001010; // -0.96128
        11'b11001011100 : out <= 16'sb11111111_00001011; // -0.96043
        11'b11001011101 : out <= 16'sb11111111_00001011; // -0.95957
        11'b11001011110 : out <= 16'sb11111111_00001011; // -0.95870
        11'b11001011111 : out <= 16'sb11111111_00001011; // -0.95783
        11'b11001100000 : out <= 16'sb11111111_00001100; // -0.95694
        11'b11001100001 : out <= 16'sb11111111_00001100; // -0.95605
        11'b11001100010 : out <= 16'sb11111111_00001100; // -0.95514
        11'b11001100011 : out <= 16'sb11111111_00001100; // -0.95423
        11'b11001100100 : out <= 16'sb11111111_00001100; // -0.95331
        11'b11001100101 : out <= 16'sb11111111_00001101; // -0.95238
        11'b11001100110 : out <= 16'sb11111111_00001101; // -0.95144
        11'b11001100111 : out <= 16'sb11111111_00001101; // -0.95049
        11'b11001101000 : out <= 16'sb11111111_00001101; // -0.94953
        11'b11001101001 : out <= 16'sb11111111_00001110; // -0.94856
        11'b11001101010 : out <= 16'sb11111111_00001110; // -0.94759
        11'b11001101011 : out <= 16'sb11111111_00001110; // -0.94660
        11'b11001101100 : out <= 16'sb11111111_00001110; // -0.94561
        11'b11001101101 : out <= 16'sb11111111_00001111; // -0.94460
        11'b11001101110 : out <= 16'sb11111111_00001111; // -0.94359
        11'b11001101111 : out <= 16'sb11111111_00001111; // -0.94257
        11'b11001110000 : out <= 16'sb11111111_00001111; // -0.94154
        11'b11001110001 : out <= 16'sb11111111_00010000; // -0.94051
        11'b11001110010 : out <= 16'sb11111111_00010000; // -0.93946
        11'b11001110011 : out <= 16'sb11111111_00010000; // -0.93840
        11'b11001110100 : out <= 16'sb11111111_00010001; // -0.93734
        11'b11001110101 : out <= 16'sb11111111_00010001; // -0.93627
        11'b11001110110 : out <= 16'sb11111111_00010001; // -0.93518
        11'b11001110111 : out <= 16'sb11111111_00010001; // -0.93409
        11'b11001111000 : out <= 16'sb11111111_00010010; // -0.93299
        11'b11001111001 : out <= 16'sb11111111_00010010; // -0.93188
        11'b11001111010 : out <= 16'sb11111111_00010010; // -0.93077
        11'b11001111011 : out <= 16'sb11111111_00010011; // -0.92964
        11'b11001111100 : out <= 16'sb11111111_00010011; // -0.92851
        11'b11001111101 : out <= 16'sb11111111_00010011; // -0.92736
        11'b11001111110 : out <= 16'sb11111111_00010011; // -0.92621
        11'b11001111111 : out <= 16'sb11111111_00010100; // -0.92505
        11'b11010000000 : out <= 16'sb11111111_00010100; // -0.92388
        11'b11010000001 : out <= 16'sb11111111_00010100; // -0.92270
        11'b11010000010 : out <= 16'sb11111111_00010101; // -0.92151
        11'b11010000011 : out <= 16'sb11111111_00010101; // -0.92032
        11'b11010000100 : out <= 16'sb11111111_00010101; // -0.91911
        11'b11010000101 : out <= 16'sb11111111_00010110; // -0.91790
        11'b11010000110 : out <= 16'sb11111111_00010110; // -0.91668
        11'b11010000111 : out <= 16'sb11111111_00010110; // -0.91545
        11'b11010001000 : out <= 16'sb11111111_00010110; // -0.91421
        11'b11010001001 : out <= 16'sb11111111_00010111; // -0.91296
        11'b11010001010 : out <= 16'sb11111111_00010111; // -0.91171
        11'b11010001011 : out <= 16'sb11111111_00010111; // -0.91044
        11'b11010001100 : out <= 16'sb11111111_00011000; // -0.90917
        11'b11010001101 : out <= 16'sb11111111_00011000; // -0.90789
        11'b11010001110 : out <= 16'sb11111111_00011000; // -0.90660
        11'b11010001111 : out <= 16'sb11111111_00011001; // -0.90530
        11'b11010010000 : out <= 16'sb11111111_00011001; // -0.90399
        11'b11010010001 : out <= 16'sb11111111_00011001; // -0.90267
        11'b11010010010 : out <= 16'sb11111111_00011010; // -0.90135
        11'b11010010011 : out <= 16'sb11111111_00011010; // -0.90002
        11'b11010010100 : out <= 16'sb11111111_00011010; // -0.89867
        11'b11010010101 : out <= 16'sb11111111_00011011; // -0.89732
        11'b11010010110 : out <= 16'sb11111111_00011011; // -0.89597
        11'b11010010111 : out <= 16'sb11111111_00011011; // -0.89460
        11'b11010011000 : out <= 16'sb11111111_00011100; // -0.89322
        11'b11010011001 : out <= 16'sb11111111_00011100; // -0.89184
        11'b11010011010 : out <= 16'sb11111111_00011101; // -0.89045
        11'b11010011011 : out <= 16'sb11111111_00011101; // -0.88905
        11'b11010011100 : out <= 16'sb11111111_00011101; // -0.88764
        11'b11010011101 : out <= 16'sb11111111_00011110; // -0.88622
        11'b11010011110 : out <= 16'sb11111111_00011110; // -0.88480
        11'b11010011111 : out <= 16'sb11111111_00011110; // -0.88336
        11'b11010100000 : out <= 16'sb11111111_00011111; // -0.88192
        11'b11010100001 : out <= 16'sb11111111_00011111; // -0.88047
        11'b11010100010 : out <= 16'sb11111111_00011111; // -0.87901
        11'b11010100011 : out <= 16'sb11111111_00100000; // -0.87755
        11'b11010100100 : out <= 16'sb11111111_00100000; // -0.87607
        11'b11010100101 : out <= 16'sb11111111_00100001; // -0.87459
        11'b11010100110 : out <= 16'sb11111111_00100001; // -0.87309
        11'b11010100111 : out <= 16'sb11111111_00100001; // -0.87160
        11'b11010101000 : out <= 16'sb11111111_00100010; // -0.87009
        11'b11010101001 : out <= 16'sb11111111_00100010; // -0.86857
        11'b11010101010 : out <= 16'sb11111111_00100011; // -0.86705
        11'b11010101011 : out <= 16'sb11111111_00100011; // -0.86551
        11'b11010101100 : out <= 16'sb11111111_00100011; // -0.86397
        11'b11010101101 : out <= 16'sb11111111_00100100; // -0.86242
        11'b11010101110 : out <= 16'sb11111111_00100100; // -0.86087
        11'b11010101111 : out <= 16'sb11111111_00100101; // -0.85930
        11'b11010110000 : out <= 16'sb11111111_00100101; // -0.85773
        11'b11010110001 : out <= 16'sb11111111_00100101; // -0.85615
        11'b11010110010 : out <= 16'sb11111111_00100110; // -0.85456
        11'b11010110011 : out <= 16'sb11111111_00100110; // -0.85296
        11'b11010110100 : out <= 16'sb11111111_00100111; // -0.85136
        11'b11010110101 : out <= 16'sb11111111_00100111; // -0.84974
        11'b11010110110 : out <= 16'sb11111111_00100111; // -0.84812
        11'b11010110111 : out <= 16'sb11111111_00101000; // -0.84649
        11'b11010111000 : out <= 16'sb11111111_00101000; // -0.84485
        11'b11010111001 : out <= 16'sb11111111_00101001; // -0.84321
        11'b11010111010 : out <= 16'sb11111111_00101001; // -0.84155
        11'b11010111011 : out <= 16'sb11111111_00101001; // -0.83989
        11'b11010111100 : out <= 16'sb11111111_00101010; // -0.83822
        11'b11010111101 : out <= 16'sb11111111_00101010; // -0.83655
        11'b11010111110 : out <= 16'sb11111111_00101011; // -0.83486
        11'b11010111111 : out <= 16'sb11111111_00101011; // -0.83317
        11'b11011000000 : out <= 16'sb11111111_00101100; // -0.83147
        11'b11011000001 : out <= 16'sb11111111_00101100; // -0.82976
        11'b11011000010 : out <= 16'sb11111111_00101101; // -0.82805
        11'b11011000011 : out <= 16'sb11111111_00101101; // -0.82632
        11'b11011000100 : out <= 16'sb11111111_00101101; // -0.82459
        11'b11011000101 : out <= 16'sb11111111_00101110; // -0.82285
        11'b11011000110 : out <= 16'sb11111111_00101110; // -0.82110
        11'b11011000111 : out <= 16'sb11111111_00101111; // -0.81935
        11'b11011001000 : out <= 16'sb11111111_00101111; // -0.81758
        11'b11011001001 : out <= 16'sb11111111_00110000; // -0.81581
        11'b11011001010 : out <= 16'sb11111111_00110000; // -0.81404
        11'b11011001011 : out <= 16'sb11111111_00110001; // -0.81225
        11'b11011001100 : out <= 16'sb11111111_00110001; // -0.81046
        11'b11011001101 : out <= 16'sb11111111_00110001; // -0.80866
        11'b11011001110 : out <= 16'sb11111111_00110010; // -0.80685
        11'b11011001111 : out <= 16'sb11111111_00110010; // -0.80503
        11'b11011010000 : out <= 16'sb11111111_00110011; // -0.80321
        11'b11011010001 : out <= 16'sb11111111_00110011; // -0.80138
        11'b11011010010 : out <= 16'sb11111111_00110100; // -0.79954
        11'b11011010011 : out <= 16'sb11111111_00110100; // -0.79769
        11'b11011010100 : out <= 16'sb11111111_00110101; // -0.79584
        11'b11011010101 : out <= 16'sb11111111_00110101; // -0.79398
        11'b11011010110 : out <= 16'sb11111111_00110110; // -0.79211
        11'b11011010111 : out <= 16'sb11111111_00110110; // -0.79023
        11'b11011011000 : out <= 16'sb11111111_00110111; // -0.78835
        11'b11011011001 : out <= 16'sb11111111_00110111; // -0.78646
        11'b11011011010 : out <= 16'sb11111111_00111000; // -0.78456
        11'b11011011011 : out <= 16'sb11111111_00111000; // -0.78265
        11'b11011011100 : out <= 16'sb11111111_00111001; // -0.78074
        11'b11011011101 : out <= 16'sb11111111_00111001; // -0.77882
        11'b11011011110 : out <= 16'sb11111111_00111010; // -0.77689
        11'b11011011111 : out <= 16'sb11111111_00111010; // -0.77495
        11'b11011100000 : out <= 16'sb11111111_00111011; // -0.77301
        11'b11011100001 : out <= 16'sb11111111_00111011; // -0.77106
        11'b11011100010 : out <= 16'sb11111111_00111100; // -0.76910
        11'b11011100011 : out <= 16'sb11111111_00111100; // -0.76714
        11'b11011100100 : out <= 16'sb11111111_00111101; // -0.76517
        11'b11011100101 : out <= 16'sb11111111_00111101; // -0.76319
        11'b11011100110 : out <= 16'sb11111111_00111110; // -0.76120
        11'b11011100111 : out <= 16'sb11111111_00111110; // -0.75921
        11'b11011101000 : out <= 16'sb11111111_00111111; // -0.75721
        11'b11011101001 : out <= 16'sb11111111_00111111; // -0.75520
        11'b11011101010 : out <= 16'sb11111111_01000000; // -0.75319
        11'b11011101011 : out <= 16'sb11111111_01000000; // -0.75117
        11'b11011101100 : out <= 16'sb11111111_01000001; // -0.74914
        11'b11011101101 : out <= 16'sb11111111_01000001; // -0.74710
        11'b11011101110 : out <= 16'sb11111111_01000010; // -0.74506
        11'b11011101111 : out <= 16'sb11111111_01000010; // -0.74301
        11'b11011110000 : out <= 16'sb11111111_01000011; // -0.74095
        11'b11011110001 : out <= 16'sb11111111_01000011; // -0.73889
        11'b11011110010 : out <= 16'sb11111111_01000100; // -0.73682
        11'b11011110011 : out <= 16'sb11111111_01000100; // -0.73474
        11'b11011110100 : out <= 16'sb11111111_01000101; // -0.73265
        11'b11011110101 : out <= 16'sb11111111_01000101; // -0.73056
        11'b11011110110 : out <= 16'sb11111111_01000110; // -0.72846
        11'b11011110111 : out <= 16'sb11111111_01000111; // -0.72636
        11'b11011111000 : out <= 16'sb11111111_01000111; // -0.72425
        11'b11011111001 : out <= 16'sb11111111_01001000; // -0.72213
        11'b11011111010 : out <= 16'sb11111111_01001000; // -0.72000
        11'b11011111011 : out <= 16'sb11111111_01001001; // -0.71787
        11'b11011111100 : out <= 16'sb11111111_01001001; // -0.71573
        11'b11011111101 : out <= 16'sb11111111_01001010; // -0.71358
        11'b11011111110 : out <= 16'sb11111111_01001010; // -0.71143
        11'b11011111111 : out <= 16'sb11111111_01001011; // -0.70927
        11'b11100000000 : out <= 16'sb11111111_01001011; // -0.70711
        11'b11100000001 : out <= 16'sb11111111_01001100; // -0.70493
        11'b11100000010 : out <= 16'sb11111111_01001101; // -0.70275
        11'b11100000011 : out <= 16'sb11111111_01001101; // -0.70057
        11'b11100000100 : out <= 16'sb11111111_01001110; // -0.69838
        11'b11100000101 : out <= 16'sb11111111_01001110; // -0.69618
        11'b11100000110 : out <= 16'sb11111111_01001111; // -0.69397
        11'b11100000111 : out <= 16'sb11111111_01001111; // -0.69176
        11'b11100001000 : out <= 16'sb11111111_01010000; // -0.68954
        11'b11100001001 : out <= 16'sb11111111_01010001; // -0.68732
        11'b11100001010 : out <= 16'sb11111111_01010001; // -0.68508
        11'b11100001011 : out <= 16'sb11111111_01010010; // -0.68285
        11'b11100001100 : out <= 16'sb11111111_01010010; // -0.68060
        11'b11100001101 : out <= 16'sb11111111_01010011; // -0.67835
        11'b11100001110 : out <= 16'sb11111111_01010011; // -0.67609
        11'b11100001111 : out <= 16'sb11111111_01010100; // -0.67383
        11'b11100010000 : out <= 16'sb11111111_01010101; // -0.67156
        11'b11100010001 : out <= 16'sb11111111_01010101; // -0.66928
        11'b11100010010 : out <= 16'sb11111111_01010110; // -0.66700
        11'b11100010011 : out <= 16'sb11111111_01010110; // -0.66471
        11'b11100010100 : out <= 16'sb11111111_01010111; // -0.66242
        11'b11100010101 : out <= 16'sb11111111_01011000; // -0.66011
        11'b11100010110 : out <= 16'sb11111111_01011000; // -0.65781
        11'b11100010111 : out <= 16'sb11111111_01011001; // -0.65549
        11'b11100011000 : out <= 16'sb11111111_01011001; // -0.65317
        11'b11100011001 : out <= 16'sb11111111_01011010; // -0.65085
        11'b11100011010 : out <= 16'sb11111111_01011010; // -0.64851
        11'b11100011011 : out <= 16'sb11111111_01011011; // -0.64618
        11'b11100011100 : out <= 16'sb11111111_01011100; // -0.64383
        11'b11100011101 : out <= 16'sb11111111_01011100; // -0.64148
        11'b11100011110 : out <= 16'sb11111111_01011101; // -0.63912
        11'b11100011111 : out <= 16'sb11111111_01011101; // -0.63676
        11'b11100100000 : out <= 16'sb11111111_01011110; // -0.63439
        11'b11100100001 : out <= 16'sb11111111_01011111; // -0.63202
        11'b11100100010 : out <= 16'sb11111111_01011111; // -0.62964
        11'b11100100011 : out <= 16'sb11111111_01100000; // -0.62725
        11'b11100100100 : out <= 16'sb11111111_01100001; // -0.62486
        11'b11100100101 : out <= 16'sb11111111_01100001; // -0.62246
        11'b11100100110 : out <= 16'sb11111111_01100010; // -0.62006
        11'b11100100111 : out <= 16'sb11111111_01100010; // -0.61765
        11'b11100101000 : out <= 16'sb11111111_01100011; // -0.61523
        11'b11100101001 : out <= 16'sb11111111_01100100; // -0.61281
        11'b11100101010 : out <= 16'sb11111111_01100100; // -0.61038
        11'b11100101011 : out <= 16'sb11111111_01100101; // -0.60795
        11'b11100101100 : out <= 16'sb11111111_01100101; // -0.60551
        11'b11100101101 : out <= 16'sb11111111_01100110; // -0.60307
        11'b11100101110 : out <= 16'sb11111111_01100111; // -0.60062
        11'b11100101111 : out <= 16'sb11111111_01100111; // -0.59816
        11'b11100110000 : out <= 16'sb11111111_01101000; // -0.59570
        11'b11100110001 : out <= 16'sb11111111_01101001; // -0.59323
        11'b11100110010 : out <= 16'sb11111111_01101001; // -0.59076
        11'b11100110011 : out <= 16'sb11111111_01101010; // -0.58828
        11'b11100110100 : out <= 16'sb11111111_01101011; // -0.58580
        11'b11100110101 : out <= 16'sb11111111_01101011; // -0.58331
        11'b11100110110 : out <= 16'sb11111111_01101100; // -0.58081
        11'b11100110111 : out <= 16'sb11111111_01101100; // -0.57831
        11'b11100111000 : out <= 16'sb11111111_01101101; // -0.57581
        11'b11100111001 : out <= 16'sb11111111_01101110; // -0.57330
        11'b11100111010 : out <= 16'sb11111111_01101110; // -0.57078
        11'b11100111011 : out <= 16'sb11111111_01101111; // -0.56826
        11'b11100111100 : out <= 16'sb11111111_01110000; // -0.56573
        11'b11100111101 : out <= 16'sb11111111_01110000; // -0.56320
        11'b11100111110 : out <= 16'sb11111111_01110001; // -0.56066
        11'b11100111111 : out <= 16'sb11111111_01110010; // -0.55812
        11'b11101000000 : out <= 16'sb11111111_01110010; // -0.55557
        11'b11101000001 : out <= 16'sb11111111_01110011; // -0.55302
        11'b11101000010 : out <= 16'sb11111111_01110100; // -0.55046
        11'b11101000011 : out <= 16'sb11111111_01110100; // -0.54789
        11'b11101000100 : out <= 16'sb11111111_01110101; // -0.54532
        11'b11101000101 : out <= 16'sb11111111_01110110; // -0.54275
        11'b11101000110 : out <= 16'sb11111111_01110110; // -0.54017
        11'b11101000111 : out <= 16'sb11111111_01110111; // -0.53759
        11'b11101001000 : out <= 16'sb11111111_01111000; // -0.53500
        11'b11101001001 : out <= 16'sb11111111_01111000; // -0.53240
        11'b11101001010 : out <= 16'sb11111111_01111001; // -0.52980
        11'b11101001011 : out <= 16'sb11111111_01111010; // -0.52720
        11'b11101001100 : out <= 16'sb11111111_01111010; // -0.52459
        11'b11101001101 : out <= 16'sb11111111_01111011; // -0.52198
        11'b11101001110 : out <= 16'sb11111111_01111100; // -0.51936
        11'b11101001111 : out <= 16'sb11111111_01111100; // -0.51673
        11'b11101010000 : out <= 16'sb11111111_01111101; // -0.51410
        11'b11101010001 : out <= 16'sb11111111_01111110; // -0.51147
        11'b11101010010 : out <= 16'sb11111111_01111110; // -0.50883
        11'b11101010011 : out <= 16'sb11111111_01111111; // -0.50619
        11'b11101010100 : out <= 16'sb11111111_10000000; // -0.50354
        11'b11101010101 : out <= 16'sb11111111_10000000; // -0.50089
        11'b11101010110 : out <= 16'sb11111111_10000001; // -0.49823
        11'b11101010111 : out <= 16'sb11111111_10000010; // -0.49557
        11'b11101011000 : out <= 16'sb11111111_10000010; // -0.49290
        11'b11101011001 : out <= 16'sb11111111_10000011; // -0.49023
        11'b11101011010 : out <= 16'sb11111111_10000100; // -0.48755
        11'b11101011011 : out <= 16'sb11111111_10000100; // -0.48487
        11'b11101011100 : out <= 16'sb11111111_10000101; // -0.48218
        11'b11101011101 : out <= 16'sb11111111_10000110; // -0.47949
        11'b11101011110 : out <= 16'sb11111111_10000110; // -0.47680
        11'b11101011111 : out <= 16'sb11111111_10000111; // -0.47410
        11'b11101100000 : out <= 16'sb11111111_10001000; // -0.47140
        11'b11101100001 : out <= 16'sb11111111_10001001; // -0.46869
        11'b11101100010 : out <= 16'sb11111111_10001001; // -0.46598
        11'b11101100011 : out <= 16'sb11111111_10001010; // -0.46326
        11'b11101100100 : out <= 16'sb11111111_10001011; // -0.46054
        11'b11101100101 : out <= 16'sb11111111_10001011; // -0.45781
        11'b11101100110 : out <= 16'sb11111111_10001100; // -0.45508
        11'b11101100111 : out <= 16'sb11111111_10001101; // -0.45235
        11'b11101101000 : out <= 16'sb11111111_10001101; // -0.44961
        11'b11101101001 : out <= 16'sb11111111_10001110; // -0.44687
        11'b11101101010 : out <= 16'sb11111111_10001111; // -0.44412
        11'b11101101011 : out <= 16'sb11111111_10010000; // -0.44137
        11'b11101101100 : out <= 16'sb11111111_10010000; // -0.43862
        11'b11101101101 : out <= 16'sb11111111_10010001; // -0.43586
        11'b11101101110 : out <= 16'sb11111111_10010010; // -0.43309
        11'b11101101111 : out <= 16'sb11111111_10010010; // -0.43033
        11'b11101110000 : out <= 16'sb11111111_10010011; // -0.42756
        11'b11101110001 : out <= 16'sb11111111_10010100; // -0.42478
        11'b11101110010 : out <= 16'sb11111111_10010100; // -0.42200
        11'b11101110011 : out <= 16'sb11111111_10010101; // -0.41922
        11'b11101110100 : out <= 16'sb11111111_10010110; // -0.41643
        11'b11101110101 : out <= 16'sb11111111_10010111; // -0.41364
        11'b11101110110 : out <= 16'sb11111111_10010111; // -0.41084
        11'b11101110111 : out <= 16'sb11111111_10011000; // -0.40804
        11'b11101111000 : out <= 16'sb11111111_10011001; // -0.40524
        11'b11101111001 : out <= 16'sb11111111_10011001; // -0.40243
        11'b11101111010 : out <= 16'sb11111111_10011010; // -0.39962
        11'b11101111011 : out <= 16'sb11111111_10011011; // -0.39681
        11'b11101111100 : out <= 16'sb11111111_10011100; // -0.39399
        11'b11101111101 : out <= 16'sb11111111_10011100; // -0.39117
        11'b11101111110 : out <= 16'sb11111111_10011101; // -0.38835
        11'b11101111111 : out <= 16'sb11111111_10011110; // -0.38552
        11'b11110000000 : out <= 16'sb11111111_10011111; // -0.38268
        11'b11110000001 : out <= 16'sb11111111_10011111; // -0.37985
        11'b11110000010 : out <= 16'sb11111111_10100000; // -0.37701
        11'b11110000011 : out <= 16'sb11111111_10100001; // -0.37416
        11'b11110000100 : out <= 16'sb11111111_10100001; // -0.37132
        11'b11110000101 : out <= 16'sb11111111_10100010; // -0.36847
        11'b11110000110 : out <= 16'sb11111111_10100011; // -0.36561
        11'b11110000111 : out <= 16'sb11111111_10100100; // -0.36276
        11'b11110001000 : out <= 16'sb11111111_10100100; // -0.35990
        11'b11110001001 : out <= 16'sb11111111_10100101; // -0.35703
        11'b11110001010 : out <= 16'sb11111111_10100110; // -0.35416
        11'b11110001011 : out <= 16'sb11111111_10100111; // -0.35129
        11'b11110001100 : out <= 16'sb11111111_10100111; // -0.34842
        11'b11110001101 : out <= 16'sb11111111_10101000; // -0.34554
        11'b11110001110 : out <= 16'sb11111111_10101001; // -0.34266
        11'b11110001111 : out <= 16'sb11111111_10101010; // -0.33978
        11'b11110010000 : out <= 16'sb11111111_10101010; // -0.33689
        11'b11110010001 : out <= 16'sb11111111_10101011; // -0.33400
        11'b11110010010 : out <= 16'sb11111111_10101100; // -0.33111
        11'b11110010011 : out <= 16'sb11111111_10101100; // -0.32821
        11'b11110010100 : out <= 16'sb11111111_10101101; // -0.32531
        11'b11110010101 : out <= 16'sb11111111_10101110; // -0.32241
        11'b11110010110 : out <= 16'sb11111111_10101111; // -0.31950
        11'b11110010111 : out <= 16'sb11111111_10101111; // -0.31659
        11'b11110011000 : out <= 16'sb11111111_10110000; // -0.31368
        11'b11110011001 : out <= 16'sb11111111_10110001; // -0.31077
        11'b11110011010 : out <= 16'sb11111111_10110010; // -0.30785
        11'b11110011011 : out <= 16'sb11111111_10110010; // -0.30493
        11'b11110011100 : out <= 16'sb11111111_10110011; // -0.30201
        11'b11110011101 : out <= 16'sb11111111_10110100; // -0.29908
        11'b11110011110 : out <= 16'sb11111111_10110101; // -0.29615
        11'b11110011111 : out <= 16'sb11111111_10110101; // -0.29322
        11'b11110100000 : out <= 16'sb11111111_10110110; // -0.29028
        11'b11110100001 : out <= 16'sb11111111_10110111; // -0.28735
        11'b11110100010 : out <= 16'sb11111111_10111000; // -0.28441
        11'b11110100011 : out <= 16'sb11111111_10111000; // -0.28146
        11'b11110100100 : out <= 16'sb11111111_10111001; // -0.27852
        11'b11110100101 : out <= 16'sb11111111_10111010; // -0.27557
        11'b11110100110 : out <= 16'sb11111111_10111011; // -0.27262
        11'b11110100111 : out <= 16'sb11111111_10111011; // -0.26967
        11'b11110101000 : out <= 16'sb11111111_10111100; // -0.26671
        11'b11110101001 : out <= 16'sb11111111_10111101; // -0.26375
        11'b11110101010 : out <= 16'sb11111111_10111110; // -0.26079
        11'b11110101011 : out <= 16'sb11111111_10111110; // -0.25783
        11'b11110101100 : out <= 16'sb11111111_10111111; // -0.25487
        11'b11110101101 : out <= 16'sb11111111_11000000; // -0.25190
        11'b11110101110 : out <= 16'sb11111111_11000001; // -0.24893
        11'b11110101111 : out <= 16'sb11111111_11000010; // -0.24596
        11'b11110110000 : out <= 16'sb11111111_11000010; // -0.24298
        11'b11110110001 : out <= 16'sb11111111_11000011; // -0.24000
        11'b11110110010 : out <= 16'sb11111111_11000100; // -0.23702
        11'b11110110011 : out <= 16'sb11111111_11000101; // -0.23404
        11'b11110110100 : out <= 16'sb11111111_11000101; // -0.23106
        11'b11110110101 : out <= 16'sb11111111_11000110; // -0.22807
        11'b11110110110 : out <= 16'sb11111111_11000111; // -0.22508
        11'b11110110111 : out <= 16'sb11111111_11001000; // -0.22209
        11'b11110111000 : out <= 16'sb11111111_11001000; // -0.21910
        11'b11110111001 : out <= 16'sb11111111_11001001; // -0.21611
        11'b11110111010 : out <= 16'sb11111111_11001010; // -0.21311
        11'b11110111011 : out <= 16'sb11111111_11001011; // -0.21011
        11'b11110111100 : out <= 16'sb11111111_11001011; // -0.20711
        11'b11110111101 : out <= 16'sb11111111_11001100; // -0.20411
        11'b11110111110 : out <= 16'sb11111111_11001101; // -0.20110
        11'b11110111111 : out <= 16'sb11111111_11001110; // -0.19810
        11'b11111000000 : out <= 16'sb11111111_11001111; // -0.19509
        11'b11111000001 : out <= 16'sb11111111_11001111; // -0.19208
        11'b11111000010 : out <= 16'sb11111111_11010000; // -0.18907
        11'b11111000011 : out <= 16'sb11111111_11010001; // -0.18606
        11'b11111000100 : out <= 16'sb11111111_11010010; // -0.18304
        11'b11111000101 : out <= 16'sb11111111_11010010; // -0.18002
        11'b11111000110 : out <= 16'sb11111111_11010011; // -0.17700
        11'b11111000111 : out <= 16'sb11111111_11010100; // -0.17398
        11'b11111001000 : out <= 16'sb11111111_11010101; // -0.17096
        11'b11111001001 : out <= 16'sb11111111_11010110; // -0.16794
        11'b11111001010 : out <= 16'sb11111111_11010110; // -0.16491
        11'b11111001011 : out <= 16'sb11111111_11010111; // -0.16189
        11'b11111001100 : out <= 16'sb11111111_11011000; // -0.15886
        11'b11111001101 : out <= 16'sb11111111_11011001; // -0.15583
        11'b11111001110 : out <= 16'sb11111111_11011001; // -0.15280
        11'b11111001111 : out <= 16'sb11111111_11011010; // -0.14976
        11'b11111010000 : out <= 16'sb11111111_11011011; // -0.14673
        11'b11111010001 : out <= 16'sb11111111_11011100; // -0.14370
        11'b11111010010 : out <= 16'sb11111111_11011100; // -0.14066
        11'b11111010011 : out <= 16'sb11111111_11011101; // -0.13762
        11'b11111010100 : out <= 16'sb11111111_11011110; // -0.13458
        11'b11111010101 : out <= 16'sb11111111_11011111; // -0.13154
        11'b11111010110 : out <= 16'sb11111111_11100000; // -0.12850
        11'b11111010111 : out <= 16'sb11111111_11100000; // -0.12545
        11'b11111011000 : out <= 16'sb11111111_11100001; // -0.12241
        11'b11111011001 : out <= 16'sb11111111_11100010; // -0.11937
        11'b11111011010 : out <= 16'sb11111111_11100011; // -0.11632
        11'b11111011011 : out <= 16'sb11111111_11100100; // -0.11327
        11'b11111011100 : out <= 16'sb11111111_11100100; // -0.11022
        11'b11111011101 : out <= 16'sb11111111_11100101; // -0.10717
        11'b11111011110 : out <= 16'sb11111111_11100110; // -0.10412
        11'b11111011111 : out <= 16'sb11111111_11100111; // -0.10107
        11'b11111100000 : out <= 16'sb11111111_11100111; // -0.09802
        11'b11111100001 : out <= 16'sb11111111_11101000; // -0.09496
        11'b11111100010 : out <= 16'sb11111111_11101001; // -0.09191
        11'b11111100011 : out <= 16'sb11111111_11101010; // -0.08885
        11'b11111100100 : out <= 16'sb11111111_11101011; // -0.08580
        11'b11111100101 : out <= 16'sb11111111_11101011; // -0.08274
        11'b11111100110 : out <= 16'sb11111111_11101100; // -0.07968
        11'b11111100111 : out <= 16'sb11111111_11101101; // -0.07662
        11'b11111101000 : out <= 16'sb11111111_11101110; // -0.07356
        11'b11111101001 : out <= 16'sb11111111_11101110; // -0.07050
        11'b11111101010 : out <= 16'sb11111111_11101111; // -0.06744
        11'b11111101011 : out <= 16'sb11111111_11110000; // -0.06438
        11'b11111101100 : out <= 16'sb11111111_11110001; // -0.06132
        11'b11111101101 : out <= 16'sb11111111_11110010; // -0.05826
        11'b11111101110 : out <= 16'sb11111111_11110010; // -0.05520
        11'b11111101111 : out <= 16'sb11111111_11110011; // -0.05213
        11'b11111110000 : out <= 16'sb11111111_11110100; // -0.04907
        11'b11111110001 : out <= 16'sb11111111_11110101; // -0.04600
        11'b11111110010 : out <= 16'sb11111111_11110110; // -0.04294
        11'b11111110011 : out <= 16'sb11111111_11110110; // -0.03987
        11'b11111110100 : out <= 16'sb11111111_11110111; // -0.03681
        11'b11111110101 : out <= 16'sb11111111_11111000; // -0.03374
        11'b11111110110 : out <= 16'sb11111111_11111001; // -0.03067
        11'b11111110111 : out <= 16'sb11111111_11111001; // -0.02761
        11'b11111111000 : out <= 16'sb11111111_11111010; // -0.02454
        11'b11111111001 : out <= 16'sb11111111_11111011; // -0.02147
        11'b11111111010 : out <= 16'sb11111111_11111100; // -0.01841
        11'b11111111011 : out <= 16'sb11111111_11111101; // -0.01534
        11'b11111111100 : out <= 16'sb11111111_11111101; // -0.01227
        11'b11111111101 : out <= 16'sb11111111_11111110; // -0.00920
        11'b11111111110 : out <= 16'sb11111111_11111111; // -0.00614
        11'b11111111111 : out <= 16'sb00000000_00000000; // -0.00307
        default : out <= 0;
    endcase
end

endmodule