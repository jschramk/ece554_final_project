module OutCache (
    input clk,
    input rst,
    input time_domain_done,
    input [15:0]audio_in,
    output [15:0]Audio_out[31:0],
    output ready_for_data,
    output done
);


endmodule