module DataMem #() ();

endmodule