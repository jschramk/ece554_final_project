module SemitoneLUT (
    input [4:0] in, // number of semitones
    output reg [15:0] out // frequency coefficient in 16-bit fixed point with 12 fraction bits
);

always @(in) begin
    case(in)
        5'b10100 : out <= 16'sb0000_011111111111; // 0.50000
        5'b10101 : out <= 16'sb0000_100001111001; // 0.52973
        5'b10110 : out <= 16'sb0000_100011111010; // 0.56123
        5'b10111 : out <= 16'sb0000_100110000011; // 0.59460
        5'b11000 : out <= 16'sb0000_101000010100; // 0.62996
        5'b11001 : out <= 16'sb0000_101010101101; // 0.66742
        5'b11010 : out <= 16'sb0000_101101010000; // 0.70711
        5'b11011 : out <= 16'sb0000_101111111100; // 0.74915
        5'b11100 : out <= 16'sb0000_110010110010; // 0.79370
        5'b11101 : out <= 16'sb0000_110101110100; // 0.84090
        5'b11110 : out <= 16'sb0000_111001000001; // 0.89090
        5'b11111 : out <= 16'sb0000_111100011010; // 0.94387
        5'b00000 : out <= 16'sb0001_000000000000; // 1.00000
        5'b00001 : out <= 16'sb0001_000011110011; // 1.05946
        5'b00010 : out <= 16'sb0001_000111110101; // 1.12246
        5'b00011 : out <= 16'sb0001_001100000110; // 1.18921
        5'b00100 : out <= 16'sb0001_010000101000; // 1.25992
        5'b00101 : out <= 16'sb0001_010101011011; // 1.33484
        5'b00110 : out <= 16'sb0001_011010100000; // 1.41421
        5'b00111 : out <= 16'sb0001_011111111001; // 1.49831
        5'b01000 : out <= 16'sb0001_100101100101; // 1.58740
        5'b01001 : out <= 16'sb0001_101011101000; // 1.68179
        5'b01010 : out <= 16'sb0001_110010000010; // 1.78180
        5'b01011 : out <= 16'sb0001_111000110100; // 1.88775
        5'b01100 : out <= 16'sb0010_000000000000; // 2.00000
        default : out <= 0;
    endcase
end

endmodule