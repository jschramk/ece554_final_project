module Fetch_tb #() ();

endmodule