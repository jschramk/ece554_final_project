module InCache (
    input clk,
    input rst,
    input FFT_ready,
    input [15:0]audio_in[31:0],
    output [15:0]freq_domain_out[2047:0],
    output ready_for_data,
    output done
);


endmodule