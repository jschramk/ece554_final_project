module MiddleCache (
    input clk,
    input rst,
    input frequency_domain_done,
    input time_domain_ready,
    input [15:0]audio_in[2047:0],
    output [15:0]audio_out,
    output ready_for_data,
    output done
);


endmodule