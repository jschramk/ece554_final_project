module Chorus (
    input clk,
    input rst,
    input en,
    input [31:0] freq_domain_in [1023:0],
    output [31:0] freq_domain_out [1023:0],
    output ready_for_data,
    output done
);


endmodule