module CPU (
    input clk,
    input rst,
    input instruction,
    input data_in,
    output data_out,
    output [2:0]freq_domain_en,
    output [2:0]time_domain_en
);


endmodule