module FetchDecodePipe #() ();

endmodule