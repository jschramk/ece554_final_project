module Memory_tb #() ();

endmodule